`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bHd8dAtEuZevg514wI81230FihTjApZisGLz1F/qBswjNjbMyz1siJ/BYE0/VKAr
idvH+z9Y7qWDivEs/6TbqnmhsxLoj274APr8KkPjS6WcbjN7lHr1Xr8d06lWBOuI
kR4uhYECKHqh0+wetq9oRbU2/hk4/mRt3d++4HnxHKjoFpj2nwYyWpZCFM3rXbn8
lE7yl2uZltiJXkv7RnhgCVLYfjRNL/jgj1qa0njFgjwqC2L9CBFtO0dtv3D7WRYq
sTCmqzbbl2wJQp3lF9X0MYV1HdHZxx5edd6SbpttPSRh9z8hV4EIIcwYCqamcVYQ
ZH/71VexX7lanW/dYcp+xJfuSpODcDi7TYV5qSAdL2+b/HVHFGC4RbhTX4Pu2UIO
RXphSPh48soMk7BlYNMABKnbeeI7SxPqKzuMyHFus7WBwIBZ4RcjxAzZdxHPeIWi
J78uDQz32IlNxoyCqTCkfBbWy9N8Cpn6LhT0UyeDTRRLVaSbk5ze7o2NrYpCUlRg
JoTvcpcWZQYK6NqkqU3ZP/kJcNkETMk5P3abG69jFPpu2psgut239e6v1T+I8w5N
Cl9fKd1VT6YT4nvuRcI+QRTYZOVn6QeazhS0zFSOZNc2IiS2zH7X/NhxUYUNCc3h
lAqGpJ+Kjj6XScQjcMHKjzYP+w8N7SpeMnp/7Y3ZPjcWYBubO/Md70XH9zS9ouVx
N9rIfaX1++JyLIZ/YxLtyYkfX3d1BmZlR0tPVNj1uQk61xqzxXZyWvczIkQ+/0Va
hiUiXofZeSgyE11CDEvpmzaFiGuvriZafOVkLGwrmTU+voRfhovN3fT+9y/J7qJY
Kc+6JU+CKWQr/DEjEB9dB7rLShoBQIBe23TkFNl3DKwseGW9ETV1+Xg7eNNgHTDG
fJE+2UFMX+f7w5lE6HAAGiBW7w93stRON9lx+2fSvzus5vW2OrGp6cfAowvdoomA
rrXA1QiNXHHS42yCieiGJ6j56X73N9hGQzY9iEV9YyjNzPNZThjC3xmUusXQ2eev
Fo2CxGsKRWDJ8owu2q0ef1l0j/KsmZY3VuzNuX6WOOAnJKbYF8JIkgU0GceuhNDS
LCG2F1cRJqAVmQaGKH5BkFMBc3T4OjOo8Imzc68l7yK5WAD1wM7L82fpA6Rc6GqD
7T/exOU+Y9jj9QUmhqXTuGquW4TMHNv4ePnQWcDckBe3abkaO+Ko+XYuNAJRlNPr
pat4pNdnNxBOxoamxOw+rA==
`protect END_PROTECTED
