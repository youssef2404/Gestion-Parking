`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MI21TirT0fzR5PVLAWE9pJb1QdzMeNBiimzOn1++NapPlxDTQ7IJj3I1tII9xUa7
3jLjO96P1j6i8dYsRC4HiJCdjLmRza92hVhNroMuXoh2Q6Uhlf3iwRjQJH8UbYbS
22Ekw+ST24N/5WemmLlCuULjfGEzluLHqWuYrDbnxhGd473y7uT6KNXBGLI9Ifei
FkHc0l4obMnONbY+3HyZVNRoGFqcwBFeUUsu2Rd7IRdGu6E54BVr6O3jylNOWKHO
Xl/j3dVRbglPuKvS7TZvgeMlSHWhyvcDd9V0QVB0hvenIHtRGM/muVkDc6IIZdyN
bTgn2lVLSPI8CryiIfMsGyWwPQwZAZviXQFVAxSOSDo3OFYvvY5yVAO/WbopOD7P
wyxPfMQYPBjV7PP3GRfC8Fmz9F15atmyaAlPuv1RnZPCNA0nkk4Gl7VXnc31MuWy
i5opK1GcgvqPoIm00wx6TM6I6DJALnXlrwAPHSeqR+JMp+KhO1QtXQXrEgQDZgCk
hfuVEFVZl+MlgjJOc14QVGBEuYngzvXmLmiKvouf1xDL2gN8V0YklrNSwI9ubI/T
bX1uj8OaLLKmkzD1uyqdXwXx4CFRLzoA62vUGK7qTTjHbwMhLixDKYXRihW+K8BD
y3Dt4tXauUAqBfvufe3rYeDN1VEyOAzGweXKGbJAoujYC88PwlU291IxcYYYNIsn
JgqyvupabuRRwDgCV7KNCjc/NmKwxmQoFXwKc36Dwe0BBUOKsgKdH5Jmkb5R+gNu
kuTxg/m/h2MoFYdbLobsFwXiPIoIcvPAjZiZA0X349g7sAIq//Phz+S0Xk4137vO
3XKT3tEOQSsDd8M+0Hj/ZSm+wmFGVXiU2lWPSI4unpPTRAKNDicoCKcHHfHQfvfC
2FxvN+Vly3a8b2hpx3OU/dOY/nZzQitUfBgUyjjrCMeAby2LJzgiiNaw3Ef6PjFG
B+Mfexdog4Rak5VwmJ2qS9GHfTq6VtWlgS/G8QStSixaL51AdP0Ef2Mvec0AwQpN
pzryOeKb7PUDZQyRvqsdab2ctsoy875ruzNIjoihn4KO2YI2Zy3jNxp94X5+CAuq
3z0PAcIE8iiIJufMnG6VPfrAJMF5wVlvJUCQAqD4vBsPixdyGNlr3O3gyePLw2Ak
k+lLCCpICppj7iAhq4hWKYRBX557+e2MrmLMOXTFO9vGHkwaeBm9qr0Djlatv1Ym
9bsC8z4qLKAgY+vNEwu62ZgvPSnFOPBN9olm+gA+QFV6UXd830GrBA9eZx0cAClh
Qk0uJp9RHbDHIusEBCA5PCujuktY9QSBR+DNwrkRM++UBBmUpGj8uabCdQiLeKOa
7LWDMt5104Vz4WTePAZwRi8X5bK0A5SyyuUAyZM16LNko3Af1Kgx1MPTF+blO3LY
C90Xgcd9R7CIwasQGcRtXtnmW2oTeKDPgbRGphVxoZ45Zn76276TlglSwWMDuRZX
iHIVN1r8PgCbaQ/gdHYmvaPjNiM+8FSfbYpQ0IZejr/QuY6V6NE176uIP8f2TEbO
pFwtw32RLlbHmZ73JE4f4eerVehiWYdJ9bpFxlAPUHw74ATz4g++/XruTB5bl7zn
j9yEkRNc9Yf8pdUQ3Msxmcaliv5TgA5DHIS/o5m3aziEA33VxydQ5qHoD3mZTnwp
kFIZrWzoWx6Ma5Dw4Zv+gW1sTrehbGLIBGiI755Pp6A/yhO2+/xt1QhKbeleRUXu
lulewoqUOl6L0ctAqEo69BOZauuE3JBDs2l5LUAn/cn0xbe23J/drwsoUmwzamfY
hUmLuoLRg4xILLOu+oJ1llqbPrGXc3wuYzlIq4r+jpjC1SSnMPi0M99KXDoTNCag
oVlV+j7EOFR7WSwAdXyvaUaccsWcarmup2ITIIFVLOqjB+XT720EyWnGeYnXl4cM
j+yy5Bc92TpqVWUPvypexMFcFVaw2QT5eyHPPY4GsvTCtXUDaXS0osC6ux5ywGYd
twvVlusmvgro0ndsQWvJNV0P6I2snbbRB88MVry66EHZFvUuv3TIfVmFaAwEA2tx
Cwvtd2BOFNYfVSlVre29a+ZPMTskThhz1pNYQFzROGVWgSovDwmP6d2zhC5z/OI0
3s7QgAQLoJaQybMpbdNIFiE3vP+BuL0GaiDWjeGnvlu1TE72ot4R2EVmmzF+ouvk
WSp6Qa8aZIB8sUAguR7vKRw6bknQd8EemB9XWENFc92BV4Td3+Ecthccznosw3KI
dEVaV6cGqoHXkh3THwYbHXIug15tfyNr4vqzVeSHr0IpF2L+8TfhrOKG3GFmjzZn
ZAI8q1CgyubMXVQhb0L9QkbZFvsKKuntbtsUgoDfajY51OtOwrXC0lju62TVBatS
D2GRf2Vvdr7hBu4K9dGMJodF06A6wcEcL1XQuOlUjWrzc0bsxsDEqiBoxnMzVcun
jD9JNQCMFQn9w+KN4UYnRiToj2fVIYE3bnOgPG828q637k9WOCIvFoJxzcYh+XQo
z4OmseAEQaUQNLLWEhT+wCm74uGfc4/UMBDU7TqbMJRarRiD23eXdlH5bMM9thqv
a4HmxuU2mcPO32a5lIY0FvigK2j0KJueceMw5tbLKWQiYo0j+NoSXOxnO04nWY27
sCVwAH0UH36t5TLS9B4RF0ct2XDbPuDp/j3eyClXD26NVnwM8XPN1sLbzJuzuGV4
FJgCiIuaAFDkN7KFTE8q8Rhmbaa8NtHrkT3yMkYJ5ch2OdTHp6NqaVotQDNOYK9q
gh4kucaH9t68mt/infr0WYaN41xpJ01zuX+YaWkYVZW85N8mQcyFcuPuJvEmKui+
hipoyAUrU12pE65hge+R9CwYknadUkCci/WzrYWeyGMRrlNMP141s7QY2txQqeFX
9sjyKFxmDATKSWxbianWoIQO5YoNpQApPA/LvRAvoLFrmicMDLM5yTM6tbBTUFuX
uZrFTmqJ/sPfizboKmZiTAQLaG4XdDtVeSRUOemB5pQTAijCUGdfo6Fx2IqO1big
5PA9r8Y91MGQAJ7xl7WbEgqLAHFjlWaAFXNvzwhMEDqpOKzlhkU9+qwTezStElt6
+NFNcYSA6fATj5IupOaz/vDFXgUzNg4raPhl5eTaItS1AoYjZ5eLP2bkCW/ftkw9
ig8V3KshN8Om1f8kKlv88vCVlm1cwL/lGbr7yKbSiWe2xuJWECytFVDXSagXANFj
DHb6g05cbZudSRrgI+/5b7r6k71rOjY0jkXBbBT/5p6fD857QjFyk0gx/FYRWdia
GclOHNSpVyO4AenX7Ye76aLFoD70huYRCpgZhQ0Hvls+Go7Dxh/5UPcb0ZNt5lpD
iHlNeB8cyT2oE4zNuOfwQ7r9l+QqWXANcatoRaWdbGWsrltNvVdj1iQx1V69NUPK
a8aFFRBPKX/zB4CDkxaQJz3RtfaEoH2AYSELPF2qNLSTx5CX76XWsqoV+VUV/19p
ohAMCAFNDmpb/pSf623Fg8ODPC7MoHut9aEmbIkTPzx8iuFz0CeXXreCoOdgATKe
2WV0XLkBc3XPgBUhRM+sqcAufFjkWXJMWMhC6YhtDXYxkBCcTONGY9ygoQtiWvrE
ajPYE90B1sWfzTHIexNd3jInC9ndmMaBhOj2ogcBmc4I08NM7u2nozCvomuFhXqq
8pkktwUUJ+amtNQoDAqfRSp01xzgDnpGIQJe1kzCspR0hicKDPKLAG6Q8elZBJYy
exy/ZqhzM+C6Fx0la85hYMn50kYzf3FIoAyhgrEkFk5ctv//MlxCQhf9j7k3ALlH
T1cJr7+ok+jPfmVtgJLYzvlKUwvtVhlkDgfgoBENHAEp0fBeapCWSgjEMIl3UOsh
R9y9AxzWKl6jqxNoUKXDXarg3vciEhjTJlrgfvqd0/oJNPXr8g5l4XCSu9X3Gi2S
25/NIOIBu67YcbujSSsr66BR+erOtq3Xtcz/EtBMVYlZaU6u38vm2Smh0uMLKIpX
ZljaqX8VNE1JJiMAwz/IxybySt+QSqce3ZTT59RNhRgB5wdtjZM3UfhbGdoVr5mY
TJJHtvw5uQiwBojb1gw3GkuiItmn4JnSFTqZ4lppaQ1bhor01toHRW8Jqja0kdM7
2czCdUwcSJGVtg7LiL0yi6SyLK3WQlE95OeIFgbLpVQf+eziNlZu8XT8GR9FlzaK
EzwNIAUZu2BkPqNx+Dbl911yF/MUrSDUJqDY3YGhkU6IdgG6qCW3jgwfFJnqwR0r
oEiX2YXcRL/ojM4b4bd+l6n8GShls0RRXjNe+p7YAkh8RmF44t9+VSXQyDuObW9r
OhWK1FGHHi5Bm7d5CQ3HMwigB6A0iG87ww2AZy8MpdVvbTFn01YiaUEq3FIXc7lp
OrHSoH8hrr2QrvH1wQfhwk7Xpzcypa6sqiNaceZwkDi0MnWkvOGwK50WZSnfFwXb
fn5mRKK7OUV82cn4LJagVCaJXOOnSlI1YfbLNAei2Obkjfhmj6Jcr8FtZRFZbcgS
o9JxHgKti1DKTR75SU/n/M8DS2pMd4J5i/bkJaEX2A8Ky/1DHZb3FOmtN1uL8qP3
ac4tUSpQ30KtDExFKVT9t505jfunlhKa/BT2DowTyHVMO5Gu0r9W99aqhmwtp4jL
z8GGACNVnulIi/6LEdDscJrAZaXCVezQZbtBA5twhT7ABi4NAr1o+mhg1Ic7glnU
uVk+veBHHB4DFthAVjWuNNIBYphAY9rK6g6SUxldnvg=
`protect END_PROTECTED
