��/  �Xt�`$�����My<~}�A��5@%z7�FH\�0��-�9EMx*1�s���v�G���n~����1cg�&Ft��ͽثc��N�i\r���y���AKK^�z��U��Z:�;��KP�B ��N��A�:����ng�DSw]u`HР_��G���<6h���LV�laD=tp8F�Xx�(c���J3v����=�I��O&��2��O�j
m�ҡ��rz�z�v	R��"�R��췰Z�ʁ�����,�>�����P��$�Y��B}�R�w�Y�["3̊���e�Hʩ�D�$���s2�l*���)f�|}3���K�q s�])a�'�<7�������0ꐿ�	�O���K�"BH8>�?�ψ��ޥ���Hd�I-�m3v	G�W=U5}��JMi=���KR5��꯼p	7���{����z��) ����lʉgv���:rf�m{v��9�3�B"���Ԩ����+�p-2�9ᔚ��Ao�J�T{���i8p]E�sd:�R�����Iv��t��s���}�'��bR2m,� �Kɾ帢���N%3gv�cٮy&��"\��m�ia�J���|_�������y�����]&L�]Ш["��|�
���Pk`�e�,'8M�X��|��4��g�	;N��P�D���i6�M:Ǔ�\
Է�l7�4ݫ�ZEܧ���k+;>��j�K"���1�6�G�^Z���.a������7/��C�v�~��yz�e4:�e�v����6� ������6��B�,��`[�"	"J�E�L��SYC�|rͽ��Jqa���3��5CO�M�i�f1x��g?�O�OR��xFF�⤻�j��B�f�
�kJ���&-)O�,�g���+K�h��1S��P�=2Q���w�����y,����a��&�A"~��k��<dmg�*/��1B�>c���g!4?��d,���9.m���_�H��lz�N�6N��~�	��K�6o�`����'<���9��$V��,|�0b+���t����b�!:BNGc�-{������	.����F��N>�ʐYN#�� ��
�y�%�YQ�V�d ��V��>c�G�v��<��4ۭ�n�~��,�gxK���U'�"خ��s�(�p}��{�8/N���@�X�BԨ:i�$zy�$���2����d+;��]h��P� gz�q|b�����!`^%�ΪIw����bK�2�,�ٙ���/�?w���eՀ�m1����ʧc�g�V*.��хF�B��;�%׻]7*�!r�1~��t����	`�8t`^�xk��i��g��p�3���E���T�4̫N�ƐO�y���jT��i�-��R�s;{����I�B��e���`�M�Y�g+|/R<+�>%��e��L�kӗQz�t�dz�~��kY��h�����6�	�\׏��~�s�G4s���7�	�ܝ���/
i�<�[�W��c[�e�5$ �������~M�W�\	�K�Au��7B1E�nj-���l멙�\/�3����v+j���,��rq�DZ�4��l��wdV���&�OkWW���&��k�!���қ��(W}&,%{j�Ս�@491@���X��FEU���/(��tq :�EA�N���<���[�k��3�����1&�+�<`�:�[�MFC���&�@ؐ��[U�C,s�RjĞ��Y>���zkJ��;��+
Z��~�Uvxn�Gu^Z.�<���3�Y�ƈ�����5���Oz��x ��� �D*F:�E��f0�I6ֹxz�t�����Mg��-��,KeC�f�P�u�!�!>����1�j��B�Ģ���O��-/Q$?�������ZEq�?(id�Q�0}
��^����h���D������`��Prib}\m1Ԁ$)������-�U�I���q#HE��Y��\��{�e���p��X�>��ټF|H,}�������l	�N��a���nh��я�����ޓ5�����t��E��f&�vt�&c����kA?�sr�;܂��ݣ�_�DÙ�.lfFv�)�c����¥�#����@���4��&(s��Xc��v��M&&�e�6�Bu.̩q{GC�հ,)����M��R%Iqcz��r�u3��::���d��)�SL��5����)S�cb��^Z����6B���y�Ȍ�L*��(^�%�����j��_���̥��ڃQj7G��h�g��_?��HD��{�/���L�*t�Z��.��%�_�&�[,>�k����������N۱쏃��"�*9wm]6�Zp���û�w!�nT��fZ�Ե�K��b���p�}���ew���[e XY��Z��r���G�(���wD� ���/�ƨ��:Jb�\LL��O�*Y2��umO{��X>u�)�"qc��� Xn�MT{@�=Qk�!��7�>ѫ,��2��ͬ�y����@�m.z��zv	:��Ǆ��A+����Q��6Z���צX���������V�|�'�7�*M�,��"��km�$��~P�rz��o���� X�v0�5� E����S����Mj��'3���W��������̠�,��?�v����5�6�h'���"�3+¶虢�����(���Mf��7f!�`�LAi���t\�oD���C87N\�GӄVDR>��D�b��|�8OaY��Q�������K��#��2ϑ1�>"㈴J�~��PA��Aj��|ԌW:�t�v�2�=�_�Z��I<�^�h9�,
EO+����*���1�o)~��X��s�3g�5��D<N�ޙ@����s}��ǩ��s��B�޵Z1��[���q2q�V�:���h�r�j���.��P}�0�T�|�ݿfڢ�5�r�c��0���,8�w�1`sٶ�E,�غ>�����%�����,��s�4�N=�M@��o��"��� GП�EV��o�b�<'�Xxfe�����qދ�xU>DVB� �Xe1�w~�g"s��W��R�;b<�<����K	3���P�wQ��U��	#�ӣ��FJ�p�g�W`{vD�Й��{�_��]~lh�Z�X���I����m������1�~ǒ�VT���!��Y�uHNX��[��k���L�m��t�֕>���Kz��(���ئ��6��h:T��S���`�uyhi@x
��9�� Ý��q���2��*����d��=q�L�Ī�M���� b���I�j���K.6_�Bq -jo���.~�u?��A���H�S�{�W�?X�Vg�sl��89��� ���:�4m����ѮW���㹉�IG/��:W=j2�2{k$3'+]{N�|G}�ȿV�>k��c1p|;�W=��8}�r��Α^�8?�A�1�RK���W����(z��Q��d��H$��과9�O��aU�x��v�q�ږ�HIh��Ƹ24w����$�貤��V\�;a�^x	(���:�Eo���e�����q�Kk1�I%ֳh�eԐ�Q�]�8!cg6�o2��k�#8�51=�Gc�\�ց�9�� �������,[]��Ta��l�߷�B<-$a�f�od� �ODT>�����^�B�gg� ���Z'�f��<?I��n!?n��*dy5j/H����ErV��M~Y����O�4���s���#��,��Ъ�R���eu�w���aƋ�Ւ�:�%2w��@~��^��|������ڕ0Y���0�lZ�JY9�b��G��m�a��GM~�a���0�#L���QO=��WP"8Ũyq��|uZ��ŝÖ u�5U��� ^w]>��"��IWῧ�M�/OM�d����6��E"*���� k����q!/����(�|�K{?Ƞ1,�y˹$)�|��
c���C�;1���[��eT�)N�MSb�i�񢻩�A��!�*�\0�/dG�<��F4<��RZnZV|������ޛ���ޡE��\��h]���R�=mv*m����QD�v>��;���X\�"��7ׁ�5 ����鯬s��"?Bp�]�����Ї�z8*��ւ���]}��y��Kh����qy�Ca��7�U�h~m�C�Kx�jR�"�KzL˭kV�Ǒ;�/��	6Q�'EJg�1B+L ѯ��{�¯#&|:�GO�si�+a_�\�]��#L=X�V���H������� ]	���iJ�Me�H�`����^yQ����=�e^"I�ef��dT���D�4�~O�`��2��`ōBԊ�Tש�%`���n�|�xZ ��a����=�`x�:0ݠOk�Gk��h�B�i�4��Q���ѿ;�w۲B�/aU9�WU��� yz|ւ���MbtR�9��̾��L5��t���K*��Ę������J��h3i�\�5,�X���m��T��L��)LI���(/`y�k��I�ͳ�PV��vd�'b����P���ɋ�6Q7.KsK����3y�A��p�rd��`kj��7b7�eG�L��d�� 5��_�c��ݛ��J�sp>�6�̘��<���)�l'.Ӣt:.=��9�!��{���}e���of��,j�,��gvϬ\��3A/8m��X��K����!��a�}9^0�P#����]b��&G]�(��6;�9i}bh�X���t���Rb=�n%֫��uY�7@p��=#�d-Y��}!���s8oF���|���q�W���o�M�}��CJВ�溫}�1��H�x2�~m��ac+�o��:R���6�Ӣܦ)u�H��t��AߟW�@�C����]2��v�ķ��xR��$�[�<�%����۰$)���6��A�+`N�<P�[�sۧ���Y�褧`���̧���7�4�ƌ��Rskt�1�]q4?��z�<�G���S�����o0����Kۆ��B���������}3}��d#�e��3��I��}u��:���g��Qc��c��
S�#�Ղ�Dx2�1Eb�ɕ���[��qg�#=1�W�`�	Z��bj��0�4�����I}�T�$U��-?����[����c�� v^�b�eH���� /S3�q��#�`�|R��8'��Z�E
OhC2�s2�o��c��1�ݻ���N��� ���uq�GN��<*u�����n��@�&bҙ'?@����k�&$����lf�f��21lm�����úC5�Ph$Ӹ���q�=0B
���#���#.��� �\y��{�c,�<�5кU����s����,� ]�{����
G�N�+�,K�I� �O�m\������f]��i5xM�.�JU5}�jP���M� b8l4�7�r�|X�.kb�&�E``O��lOL)�p���}�滮�K6�K��l-r�kɹ���T�䒣�N�ܘ�g��?�T7�ǦW�L4�m��o���R�������$�_K�Y{�M�l�;gX��'Vl�-���̀4O.J�/����7�l��g�(Z2��|�y sx �!��Ԋ0_��t��	�8s���6g<B_���|�2	2g��Z�320&u)ʞ��q����$�)?�ì}�zP�F��@c�{�#n�Ys���a��A���!֞�d=J�_�*d�HB�"��ʷٳ�=�
���Ѣ�Q.�}��
̝��#V����":\$o�`��rq���̽V@\;Ԋц���zRK�*תw� ?�c%�,@%�;�ʂ�o��}�Qz��Պ��O[Q	[�}��,��͕b�^�ka�2����憲l�h���_�����ї	Γ�ĝУ��+a�L�M^ʜ�E�)���g��j4��o~�}�?�n�ɑ�e�ݜ?��0���)�+p������xq{S 
e�5�0%oP��,Z.Q��'�i�<D�/T��v�"aE�®���ȭ��o@��]c><TV�	��/W�
��7nSn�rB	b"�6l�3��.-'R���0`��D�h?�V���V�{,�Ǝ@8Y-��K�aےvQ���Y8�mk�o���1�����m�fT[�7'ޗyZa���G�A����%i��~t����{���0���p)Jir��V�Pa�a�l K>��?V�(��vwH��q�d/_���f�:D��ͥ�A_.��/#�r-�a:��&�&(��{Vo�
pŪ�~ҷ^��)�/p�r`5��J)]kʰ���J37����&+%�J�"��.n)^���n�2w���#����(��E�RF�6�}�b\����C���,7 �I����џ��>��2��HH=�xS�>��NRna}��Uv�>v)t+��o�����SCը��KV!��!nU!-i��s�:�>Xi_�6���S�ȥ��,�&5g�$9����� `��+�d���(��ٽ�R
2<��vR��:l�Q�{ç+��Y� UY�;�d↍��NП��G�F���M�ɤ����2��X����S��s޾}��kY��'�=�f�]���)8�|� ������9.�al�^�%�[�W�8�
C^Д�=�����R�;8�����M�YF�R��i��{��m=�o���MI�a���oR4ȧ����]��lYK^���_�7G�Zz�q�}�j�Rz�3h�=���L-�1.���<��Yv$��㻼����K��� ��r��cCJ鷩��q��X�3���zu���D�O˲��b
����R�U������o���]P� ��=~ɺ��3K�b�ʎ���~���i(\�M|*������mZ���T��C[O/S���:��F�dևkМ�&�M�d�K�"�
�����~1g�biFO�djw�	��X?ǸD�w���=_C��9��O}k6�b��gQ)�R�.O{��McփO�-���Ui4�KTRg|�9�}��ܵ�t��ٽJ�f�kWW7�κ��XF�3�8�_�����v�n�>R�A��%�aǸո�Ⱚ�0�Y-?�9\=ܲ��s�xa�"��'f�*�yQ J�.; ��J�����C&�*��G.��j�A8���R��1W�^I�l���.,�S��Z�("�ze�޾MD��D<��0i�
qx6?�*� x�2V��%�{_����1�䊞_�
!��g $9��B���e���Z��i~K�ף�)*@!�ok8l�w����EF,�6� S)�p�"���x]&�YP��� ��6��A�*��8ӡy��h"���*�i�DyR��J��[��YbCCO�>�m�Ue��"G*i�И�@8BW�,*p��s����4g�Oe���H��yh\����0�=��q�/"y�7��!.!� n�m���19g�y5*0(��P��i�650�n{����� �,ar�j��݄c[UẮ���T}�I���IY[c)5�	Q�c�K��"�[I|AoE�[e���CO�}��� v�jf��*������1�ս*�9`C9�[d1���p_��2m86���+����[-��4�뉂Oܝ:K"��~�7 �M�[|���me(�+�/�_�"�[]$�/��Y��3������i��H���kМ������=��� ���O�n���c�z4��R��k��>�/l�~C`�)m�i�`Ӕ�1>(�;�go��'�o�=Huf+��!�}�N�mٓ����q����&VlbG�.�V��홽��.�	����6x����ep5S�������+����9�	�<���
;$8�|���<���ĩL
1����r�`�i菈��t��`�� ��e7�����y@GB d��Q�mk;<[���G��'#Y)�wQ��r�Qp���b��<.��Q�j�|)������;��]p&oK84n�� �{.b�Hp<Q��Y���B<)�K��.v�(�ާA�����u�9�ƅ��],
o6|��sX���J��)BJ�S ƚlc�j�4#�KT� �S3Ь�%�QR�6�aɄ��]�A���"�a$/�Ӡ�v���r!`����h�r��
o��S֝zq�?iA�q,~7hf'ʢH�Y6zD�k��Z�WKu�ÿ�(Ю �Ag����p�N��i�gl��i]�,%o���Ĵk#J��s�ڪ��B��4f}��/`�SV��7��f7�H�kX������3�]ꮪ��Ҝ2mج��?;�D�-`��]�����eI_�����:d�>��h3��~�)�%<vB�R��=��6�z�m�F���H2|��mf@����Z*9�3J.��h_5�y�&BD�tC���)ȩ8�_~����d殑 '0��Vܑ�ү���7V� �����]_�4���)����3�1� pݏv��~��������Wü��B��H���]�Qf{
�t�_N�+����!a'C�D�վ����v-H���R�4Z6VV-:kV�\v$��z�Ÿb�0#AmVG��]�Ө[W� I>:��$W�'�=���ѹ�)M����e��C鷵Q{�b��<�+(�z�4r���C����F�>����ƚЎ�F%ђ'���a�Քz��۾v�؋�ڈ�)a�a�C2�g����[�&!4N\��)��Mge4㔮�a/��w�+#x���e�\���^J~aK��M� � ��`���.����X�`�.�����g��B� ���ɜj޳��� ��k����K�u�B]M��.��2j�x �I�%3��ҹ����HXnq��(�A���S����f�I��E
���S�"�Hc��2�H�,��R�5��n)��[���!��Vfa�a���2[�O��/�NO��q�� 2��U���Vw⢠�ZC8ͷu!�T�xC�R5��-��)��2�g����n�t��)v̝͘
�9s@�á� �`��F�Vǽ�;��G�i��ʄ�a�Ǧx�H�ʻ7\�|�C;�^�\&oͧ|"/?8a7X9YMu'�*A����L3�����uFύ���SNV�'h��L\�3"��	He��v�b���B.�y�D�:�BI�d�4Ζ�2��Q����}t�sFd��/R�L�e��Lz	�¢�=݀��1�YC��vb2���Z3�u�g@?����������a��6�����9��p��f1"^��E#��l��C~��t���
�@n�<��=P~Հ���
���,�ZP��3Y,��pK��@*��"�hf GvIuqD��Lv�@?`��>���� �u�Xb|��E���,Z��B���L��������!�Co�7R,ܥu�ULVy#Yg{5ә�LB;� Ł�>�g����DO�
�3�q�Z6�Wu�⎙B�����!��?[㲒�I�i|�� �S#�˟�v���?�)T�4��cIv�!���[��Z�K	�V�s�h$Hq���LͲ��7M,,���	�&þ��2��[�	�K&U�e�1�R�>
<��U�0Ō��U������t/�Jv��<�9i�k�.��r�)���)��%����Y��6o'�ފB9��L���,����!��tB�0pZ��AS��{)i~I���9J��l�A��E ��?G�s5bc�LpȈ]}h��^���8�at���G%i̿�J���NGp����o"�c0>�d'�[���	���F�8����&�G/�?�֌�J���xL�]��^�B���-�6�g��X-s�
��t�L�S�=�*�m�o�q�����v|
7��UCW�� ?�)O�J_�2��N"�G+7�S
z\������l�Eㆤ�����c�-��}d�=Fި�c�V�N�.32��2jM^�᫣h��`��x"�q9Ǿ��Cc9�rL]�Ѱ@��I��T�ֻ�Y�\?�i1"^�~��+x��֕�i�fx�յs���(ºKec��!� e�Pu�-�C���#R�?v�1��U���e�,���>�����{����{�CӢ�}��_-���s���~��,�r7/O��O���0���2ۚH��ژT�h�� �xʛ^��|�9�Z^9�F�H\��u/�^���xO���i5�?�}{,� �>���D!z=�ѳ���#^J�dN����R3f��`d� H�.ͮ):���Fn�3`$���{��d	��S��"P/I8C|��l_QC��Q���in�u5-`�>�O�[��2B�"�
�^�h�e�[OԆǋ����U�*�,� �p��� �21��1`Q�fe�1�����j@>$���m�0�h��!��>��ۅSm����e���n}��"Ğv�!lV.��-[x�Y��_��o�5p#{<�p�@��4�2�������d
DT'b�+W8�&�&+d?���QV�J��{�ʵ���@�ύ�t�z��T-̓C�sS�J��I��j���*��������R��L6�"�g;;'�\h���zd��� ]���rڻ��`��E��{���6����~,v:^0K��!���Sn|����� f.���"�p��]���v'��٨��ܫp�WUW��C�<�g�
�B����U�!���J�@|/F�u��{|�lE��+�*D־��;�����X�&��?��E�-Ԡ_t����-���~�+͎��VW-4��]t,�k���g�����	p��Щ]�W83�5���|M� �W�S�;��5Ba*�ؗ	a۵���U�;���'�=UYz��'1߹�����&PL �w�,7:ڥv�	�P� A �p7x��ws��$̲�µ/��Ntr���Ĺ�H��	f%�5�Go& �F�>�Ɍ�-���\I���}P�e��s���a�t�{�	��rr�6�5��<��ew��2��
��q��$���ޕ��`�*������x�t��آS���u�-uJ0�E�IƂҭC�L�s����b3M���Ma�=/[iq�Ќ��ͳ�B��T!TL�I��U������-Ȇ�����G��;s�h�SQv;ב�J�6�"BK�ͬ�$A=�%�߾C���ZH��j n�mv�{��>�,���Ol�����g��R�w&�V֖��҆��H��i���_�myVDR�2��C�D�)h��ӷ��\��N�HHY^�_^z�	��_��g������m}��}_��	2*�Tv1��Xa~蝉��q!/~���&�ܠs[�d3z�h���w�dٝ��83���mt��=c�����G�I�� ���/W�wi0uZ���b������<���m-�z�,��v����#_Ū������=,��T�U���I�����+�Gp��;��Y��Py��n�N����\���cP�!�� ~;CI����&+w
C�
�w#�%��[!_�v\�jғ����ٝ�h��
��F�.�u�غ ՞�
b����W6y�9s
 �YT�ġ,y�$�4 5��ӢK	�� �{�S�S �%�����tO ]��[�Wk�, /�sbq3��kJ��<09l�¦��*r��A��6컰ꦥq�\5����c~&�����Q5�+����͈��c�9���v�D���%�� �_�Ȟ��d��� 	XX�g���������:?ˏo)���ޥ�,p�G�(#o	�8Q�{����카�$�VnXH-��jm6ypGGTӰݿ�F��C�3��J�5��Њ`X�V�f�r��c�T3'c�5߈~����:�QӜY��6|�5;��tha3Εz�\\�*#��]��q�	�������
��Jڵ��7�Q��;Pf?`]L�{��0��Leʺ�d�;����i�`�Kg�h���R��1|��E�=�٠2��WE������۞V2k\�Jx�@���ɫ q���v�5~�K�}eV*ӑ͛Ϛdv0RZ�~�/F�
�O�П���|a�ny$+��9�H�� ��*��fC~T��#�p+��^��	H��8XsKO{�S6�;<������hg�*�ɿ�!_ڈWH�b9�����	��fd�����~��=��Тz#K ?	l��*m���F���h�5�5��x��'��.Y�U%�m�_���*�G3x��BD��$&#���^l�9�*7�5�?�!�)���|Y�&w���&2=~xW����)���gXB�i�A�� ;��׮�c��Q���
s��/�}�f�/�<�oł���-2��zS<���'{"�SI��J�Y
�Xv)x�#��c�;z�%�u@v^���Y�޵pU�c�(�()z�[�΍@�t�������P`ILÊ�"/(S���f�&==�-�;¤(��ϡs���I9��\�.,C�XT �b��0�UQK�x��p�u�E#�ez�]�LA�
��]-��'��t�Ѯg�/�lW�%���}䷕`Φ����6l�����ΠҮ_�Q��y�K����������gA�bӨ��'��7[�f�~7;�#�>=8U�b�=u{6����R�0-&8��(�୸E�02�cq&��qn���Hg(*MT鄼������z&ޮ,�p���.�L�����˜���/��C��ݗ-�����	�ǚa�@�����5�.4�� -z�"���23J��v!-&��;z�cL�_�^�BW0��
f�������Þ.����,�>-��6)O�V�X�M"Hi���������_�Z���|k���ᅓp�j����(_��D3E�it �j�Њ�?_�c\U/�r�W�ghgM\�w��>��>�? ��8%+k�Ȃ&��X�bG��.`2�&렅�p�]�COmџ�W�����D�3�:���YM�Ui������[(1=�z��v=��M���c-���[ �'�(9Ö�LB:��TTV���C6�8���e;��5�}�`/��zq��.�.�D Mp��$p��)s+cޫE�\����}�[;��#��pM�(�*�a�u�I���0�v��[�W�G��c�C�����%Y�_I��0Ԫg���)5���i��'Z�wT���c�c��h ���,Jپ�����s��!#cH{�,`�� <�s�-��N//cq���|����[�$0~۾�|e2�=�%��90�X�(؎S�i3{�JD������Q��=���T��1|^����7D+��w��ʚ���/L�9�d�Kb�� �k�����Ϋ��V�\9��f�f��{:��,T���� �����ի}L�1�i�0�ƒ�]pvH��̿��
������S��h��V�ù�l;��sv�A^�dA���F��?�'�-ݝ����(�)�}a�廠zڧ�C����y�V��[��?�u��C�z�]Wn�R���+�8<(����F�b������	~B���B ژ'��k?��٫s�&9�ly�+�l��Gp�M��5UYM�$ЌV������{n8�}�|$n�P�Z������,Z���?�N�F�E/g����/���J�e��*���~����oDk]+�n�<�6=:Hb7�BR����y�%��� �g��\�����h�&�n�u�b�4���za�P���N�{��Z����f�K����\��&����\ׄ|��Ċ������!tR�K�d�S�G+�w����J�)C.�2�Y*��7W�������_�j�k�u�${��gC��Nc]�y���u��ȴט�3#٫�6��dh>p
�îcѢ6?K�-�\�!���O��)�g=�p�h�����u��<I����_3^��D�
Yi������F�ޑ���b�YW�o7�'l��U��� �<R��g���� ^����'g@W�F��2>�h��İi�����^_U���ζ����]�Jd��8׆���S& mg�����OE�I�d�I����7	1����Yb�42Y��Q��w]T��M�eG��7��7u��;���N�0�	��:HF�^���IO�=k���W��;/��c����]o��g��%��;�ץ��k_��H@9��S�h�`Ұۥ�(e�BM��&�XN��E��:_�9���J�v?�w��ó�%u@^�S7�1�P�`\ך�P�{�������u0�a\���+[J�p��9wAm�-�N9�*��B�K!�U-jdו�,t:�Ɵ��Bg���}��@)���t1X���џ�8%�=�]0=n�~� �$�n�
`�����a����n)$�?�N�i7�"�-;�\ {�z�c5,~|�
Y�t2	�k�iw�|)b��h�N#5�Mn�ֻ��$��o�`JN�9���Ъ��n����bL36+qa�F���y_��.�c��6��c����'�sJ>e1�8Sv��w��R�>VSH�na��-�$l�D��V3L��^�J�ۓr�<\�Ǥ�	�>Q�)_�~�s=z%Q`)c��ԗ�s6�.��\���R��/gߜ���*������Aރ��|Wq)H7�-_�JY���.�v�>|�{�㗞��#�y���AY69о�ONzrv{=��e}�0v���ыtji��wfd�)>�Ǚ����uK��7��I�
��*����s�6�5��R�|O�w�"�
��T(�����&�<� m@Rw8�
8��U�G�ʲ�t��9W-D��2�(�c3IÈ�����0L�^C�������[xP��-�,h�s_�,����r %��,��i?��UC�� W�[Q���}��w�jy�*Ϩ��<��$f��HVzN�-�Ju�	��!D(�Y�4o���,
v��U�7b�$C4�K�R��Q�7]a^	z�Nlu$/��J�����cpaӮe#=��Þ��,쟭,�����\s쮪Q���Fo��Q7��M�V��_����oSbӳ.�����TH..
�5�L.w۲+Cz��_c��wlHTl�M+fv���{峘�4��ᴑ*��$˴R���������{q�J����R�ߞ�I���[6��a=�Cv��<���� �rwPg�4{�Q9E� 5����roDIY�ִ�M~�����/�*� �ر%���Α�|�45�(�ԩ/V���AK�-�<�"!�|�8�@XP�6`V�{��R%zA��*P:
���B����.P�/Tτ�1�1$Q�����UH[�� �T.�JߏL�m��}pK�8?�%�*��$m��H�'����jO�_��uUA�x �k�F?������N�Hި���r��ӑ�c:Aq��a�B�?��ؚ'��}�B
�'/��@+/�l�1Ugi�߉���ּx�y�d����/,����`��V������]�+K =_:G��)�y@븊r5љhY��T��t�|pP� ���Iv7N=.G���씈�	�^|����/�|-�A�N�j�������,��3���P�~`��q^Oo+�o�|^:���־��xN�B̆�tw�?���:�"�1"�I�M)`V�|丁L��_�?����Y�{jՍ�
��=D�vꄪ(v(c�>�¡�0�E�r2�����ū����S�4������?�mǡ���h�![��ؠ�F�O��
��Qk��ʳ5s�M)c�Uj�*�U<�7X��Z�L2�<ޏMb/��� �X�����׻�G4�,�����vjr>���b�w�۹�_��h���Ţy��3>���oWT�)1%�]�Dג�r��.lycu���Dz� �d����QE�C_�hhdI�*������RR6�`D�2�x�+#I�z՚�_5"�
�F"�=H�;<��K����D�������²~nGy���;~�d�Ǔ/�^����چ���	G� [V-����2<v�q`tC�D�N���)�w��K�i�g���8e^�����H��	��<�#���W2*�zb��=R���u��]�!	IBLT�F~���m���q�ځn)����Y��&u;S�`7LM�zJ{��aK
���Z�QI� C�{��(ּVH3���%���Q �i{�xA��$�h�R��* �5j=���j/��z�+���*��uϯq#�,��5U}��['�gciƺ��^�I��L��Z��	�����e��UY��"��"�A��-G�$i�����A|�w_�z����	o�N�����x��_�n�"��4�m֯��רb�������˃z�|�XkO�u��A��H�N,-��I8A|�&�r|�:y��I!tr���^Oۇ����b���L��5�� v��w��5g�w?��y2eT!�4-w��$$É����$𡅛O���A7��i*��)�����p�`ͼ���= �gxH�����1H
T���iJ���L�>�b|'u�9��꿻\�;�V�?��ߟK$�ʚ�1:������􌃍�a;���D%���5�PQ[W��re)��|O{sƔ�ӎ�%�����Cɻ���Yt��8}���i�q-���0�xd�V���ٌ44 닱9!Z�+�wX��~�P����ӱrx�d\��o5�c�,���Z�*2ss�u���´uV;���~��(Ud�@�H��-sD�]��K5"gaw$��'�Po�����N�a� d�f���g�O%�lcW�xv5����}!�x�Y�n��2x�ƺg��b��-Y�Nr��e�S��.���	�!���}�k�b���g�E	���!7�Z�����O�1Э����s�����s5�F3M?�q�K��9?�/�/�]��v(&^�6ɡK8:�D�7��&[�P)���xjܡ\�#/�n}[%�g���*ůV�'3���I�o��/2M��2Ԧ�FG�����I�F�NΌ `��/9�U<��T�ۙ�և���{�j�7U�*Z����8�8�m�]��W)4�5��	�Q
Al~YRA�O�f��cW�m]«W�(�i�I������m��\�m��&�]�qbtz�`����:��I#���W�Fm[׈nʄH��=X�h���+;���g=�y�>qRQ��4�ؓ�ǸYhMҵce�Q\���y���R��Ka���p��ɇ����U��yO����v?6��,�\��4K�9~���P��+��!���eF�&s���ZU�5w<7W8g��E�\.@����S��rC��@p�o�w�a^����hx��gd���wЌؽ��2�m�/@F�TTtpU���ܟ�����@���d+x$fw�9���uc|7��b�y�D���@:�1��+~�����6!F:#�����EDa$,�7W�[�Ln�3��<�&��K��+�O~����#�/�Ē�Vy�������{���@)�I֔Ϋ���SQ��Q6���|1i��g�n	I����3�1b�F5�����L(:��+G�@ʺuo~yQ:�OR�N��0��m[&	����SQ8C���a�\��b�����a�ߡ�)F5EΣ)�kp�'�O��r�Z�/r�8�:p{q��c�F��t7�=j'�B��ڍ��,�D�
V ��[i�� � �\�B�����_y.5l�_��b m�)���;f�C�(�����RF{���g���#�C���������?k�h[�^��ݯ'K� o�q `��o#y�F˔��_W����*��Cy?(%��}���m�~����� ��ۭ҆������ĂH���[��j9/S��*����K(��F�B�v��g9��_��q��Z��
ti��	Ȼ|<�(�i��)��x(���]/-Oyʤ!T� ݁�h����A�6#Ð���~�81���㰼*��Q��M�C�U���=������+q����zh0�������O���	���C�r��Be�Nڀ����+/x�IHL��@�K�7��}�1,��
��V����e����r��� �Ic�C��#��3m��{��\1wn�)�!�9���ӤYڢ��
B�N󱜅�l*V{����<��~� G߇S7�q]Uº�+hX��:��Eu��D�7.�W�!|y�bb�?� ̼���OЋ����3ʤ>�{@��G-���A��-�f�^Yri��6@��m7�05Tz�k���ϯ-�
;�u���T���	�m(�U<T�y������~t�����)�Oa��broj/���^^���7.*��>�G]ц)��Gwǌ�si�q�r�j�s�R\Xp�%F��C�~#�'˖kk{6�S3kχ��6����B��dw�m������7���G�	�>K��p�'�l��,B��4�R�_�����)7�����T�Bb��xW-�e^��˦ -ѳ��ik����}?}Xx��Gx	C��TI8�;sK�
��0<`@E9ݢE� �3�e.�9>DS�ko\�p��c�[��Z,&
Ѱa���/�.��x��!-�2�Ĳ�(�	>�&t�`�\O���u�$2�!�S`�YP�S?A�b���}֙������B���,�	���J�Ё{[����k��̋�vB�9P�ހ,��:����T�5/(
bsW��=�"e�N7�e�CjLL�
2Xa�[f(�����������, �4�e�3H��JY���IG��=�f���]��[�	��3��d���!r��E���L/Zn�s�����XCa������'��H#5S��鈟w�Y�[���D�>�_ԨC\*���Mr��'���1^ʢ�x3�S JЩ4tx謜��\��4��c2�/�$���(@��,�h �G6�a��4�.4R�I�_iĝ�f�����Vȹ ��u�l�ힼ�a/��[���&J$i�ƒ�fm/&�Uu��?-�y�f�U���A��Ű�d}?�px{j��E���m�x�0G����R$�:7�S\7��k$'4-��x�X�B]L��l�vre���4(��5N}�l��#�^ʴ2Jˢ�i��4�8��z7*�g�"���&�p�P�U�EJ�rf;�](���టh9?��<#B̲Nn�Gcc_8?�pf36�G�l���J(婅���9?�D����� �-��L*gP���RH�XI@�Ǆ]˼a�E�m��ϣ�eb=r-���ʪ~C�?�j����I!��N���������}\���A��g̎CnO_v��p8��0���S�}p��{�n#�d>�bOǣ2/�3�[��h�~�3~�*b�d9�7eqM:|��=}ǖH��FZ�*Z��u�b� ;
s9����K-�௙ËX$*|rS9���,�Kv����C�o�i��{b��������9�k��op������6�!L���N+���!�e��,���������F1�x/q��)���$j�Z���|)k(m7]XĔa�;��[ji$���+ҝ'��|�\G�B�f��e��/f1	_�/�'�%�0ap.Ut$��ϫ��򱞼�L��X�f\���Sbg�OR֪��NM�c�W#�r��'� ����������t
[ׯ��A�z���k��o�#���Λ� R�ix=N|}�j��E��i�(���?o��׍�-�1?�Za��ex�ζ ѣ�ivi�$�+�r�iv�s�^'j��̆o{�V���`[u��S��V��	�C�B��EhQ��?|�S����0+w?�܆#��`^�9�V����=��\-���H�!Ӊ����_�q��G�L�{�ڻ�M��z�X�l��fl��T1�*����졺�'o��h�EN�7���u,�4Ŏ���\���e�4I�'�#��͍P��4�	��2l����8��-�ªȹ�e׳��Z��װ�)�GI���g�Ŕ+�'�!)4h�J�����'�pz�yW�����J>�'�8�5X������m��I:B�%�s��@p\�$��"�|���6V۽Ra���E��Lm�qFpb��Y	��T�f1�!���kJ������"8��� f���i�+�&$��U����8~�KƯ!������l{�H1��/yD����"��i��֧��n�I���i�L��6;9gk�R��ܩ,;�u1���T�$�/�{=rAE|+�=�HQt�)6Ep�#-1�h�=�v��%�d�_.�A���dm�mk�qC�lQc׸�4^/n8�t�IN�Jc����J��H[��FU��l�A.	���;M�)�x��cjJ���_�հ?�� O�TJՑ@$	Q�B�q�B�@*~��|s��S���&���lD�ڞ糅:X������es[l��	rP!M�mr5�[��8��8��,�s�F,�\ �h���	�3����?�եen:�r&�JQ�ЄO	��p�<t&�j#>���mַkH�2@��iQTk]j���YN�	����_IV��ԓ����	F�m�z�9��*��'2ӱE�C�'�qq�ߨ�1˩�[���o��(���(�cM����ʘ�q�0aɜ�|�m��3�
�vwA�)�d�!s�y^7��`�?Ač��r�rmZZl�*� ��n���h*LE<���P�խ�|g�[>���؊�m��q �"�b��ɯp!��ӾbX���(OS�@v*�>�#,�P���^<����^��6��R���,�QOڀpD�m��d�gR��/^��/��W��J���̢�пb�9�G%�� # �V�B*f�v��"�CwR�&�B=���5�4����f�=����/����-L� 꾄/|֏��?��$�Y��68+Ѐ�_�R�U�I��1�@ź�cP�@�S�A77�>�C�
���	�z�=�%�\B�.��~��ÌF��A\J%���z�IݻA�e��,��-��3���n��xo��K!�PI���㾃O"��O|�����j{�N {�L�Sύ��Y��q��|9r^���.-'�WY����z�n}H��,�]�r���9��� 8�q-�Dx�w�qP"0/�;ǰӡƝf�)��<�'v� y���%�]�L:Όr1leaK��(�2$YH�0�W�'���W�����.8b��L�ف!+.)ٗ��q�$�=�>�\���j��*Ý���Z_?Z���&PXy��S�s��w��}Q�:���u�k*,}��.�j�	�'�b����a  ���Q�^ѳ�<�q��4D���B�㑦Ҋ��ۀ�A�u���㕜f�,F��Z=ժ�:�p����F���zZ�E�+��}���f.��z~C���y��
q���H�EZ1���]����n;��H�GL4P��}m��C�ɵ�I;�����k˘7ßAWdX|������3w�4�(&�F�j��j�?��s��<H��T��舅�gwI�O��>}���~2�����9�<2��T�����m���5��[$��ߵ�Ս�dk�7���r��Sɤ��|��J�3����G��ӏ]��,�l�f�v+�� S"W��ӓ�(`$c6��.�$���ɛm ��+N���d���U]'�����rl�J�۪�U�:�����En�}�0��d])h��	;�G+�Np97a����'G{!�kKW�F���6�"[�nGS!����a2b�5߂�ҙ�����رS��}����R���
�ǟ��fV���|e5
	x�ev{�u/.^{^�X���O�E$e������K;{c�=�TF�ewY�>��Bm.��n��{�Kq�xЎJF���B�׭?'�Ԙ���>��7���%�?.����������`�(�5�Y�݉�c_���f�M�9�2VrP��8��Ѓrո�5�45��Y�T�x�P�C��_�i1�]/p��(���ξn���|m��u]�A�;�BY\��O'=#EW�Y��JJo�ӿo��m�q!O�b*�Q�hK�N|&��CQ�v�l`��ӎ��1�b�P��:���D���Ve
�Qc�X���m�����p;�����Қ##|���[*�\.���gu��;�Є��3b�7��u�sY�1v���9�ʺB#^kj?̥�č}t�j��}�i��s,j�j�7"�I��̵K�Nݘ:<xr�G�:6���Aь��|��L�Sb��j>�H�N���4»���MBC�_rX�,��}�6ɧ��iie���*��f 
1ʝ4��:0�:���ٗ�e�.֋c.�#�L�EA�1d<+73��>���S�4:d����.D�eCy8rŦ�"��p\�v��E�ܛ�3D㤞�>��m���M��=D̋,c�Z��g �y�=�$J�s2������و5�hڢ#^^Ñ�%=��"��G�� ZH�=)�}ت��i�Xv�֢\�t��$����>��#�AN>ٰu�n/�'��cbU�\e�R�| ����_��[:� p�5f����R�z�D�Bt{,�zQ�%\_ܔ��M�ۘ'�@_r�GTy�S՘����t ��\�� ˾�y���i*#v
*����*����~��F=�;J�W��Tw�b�ɋ��~ȉg�	�Rt�tÖ�!����;�o+U��6�'�+A���(�1�.z�[aDS��~�a��)�z�hj`�.�V��+1�c�d��3Ev#�$�Y=6�['F��i��<C�PC$m���� -?�n��2s�`N���7��D��#@�jL���"��*Ͽ |����8"�v��V04M�-�u�����:�����K�du���"�����S�Q�DKkI��"�L���-��]vT��ܸ�a�c���`N�M��_�!�tχ��r2KR�$�I|�
��C'����b����H�����ۇ7�c�
[Ò�t(�R�����nu�fG�kA�p^�={.��a_m̲�gD(�^��TY�R)w���U|�٣�|��-$� �p�F��:]x����$�I;��dΝ�o,�W�t���>�I�e�xR���sT1Wi� '/�� �p��գ���A��_���{ȹ{�`��H�J��>Ckr��}�0���S�"�$>�;�xU�A����+�8~�`�a��|��P#l����	�Յ�v6�[�E�:9��+�<M�r3���<�pv��Ey±[sǢ2��yy�2�@�N��M���i5T��Βڃrr�m�pv����Y<�S����P�X\�v�2�qcW;ϫ��A��BgMR4�m�?O�	�?�!�я��2-��u0�jL�p�5�&ĸ��o;��r�Q+A�O3VA$� ���`'1�g�x��xg�0Bn��Ii�>�`�C[��9$�}/g~�����˚W�}{�d�%���h΅,���E�n���q:y)	PM
�c���k>�?�3ћ�����,����ř��@,�_���m��y�����e�j�B$h�C_��HA��&�Nh����X�5�`fy��O'�ڎ��SV5+��,��y��]ƕ��J͍��@��l�	oB�<K>��q@��MJ�R�����Ҥ������;B���Ӧ"k^�Ì� .��� �3 5�zC��f�̮mT��/�ǯ�߀�_�R�Y~��* �*Q�dh��U�gx��ϥ1���Ts��fڧU�Jք0���� ���o�^qS�*
I������ZV�ĉ�:h�n+�B~�����r�/���di��M�����������.y�r��D�(fn�۫v{M� �c]�Zꕂ��Mk��p���*��_�7I ���r���#û���ft �����ǚ��D��C�RE$���
�Bl.i���\� }z9�/�m^��N�J�I��Uob&q;`�`���]q���Q�8�M΂� �8��qT�Hx����1�s}�U|�sEl�{��»��}���Э��k�L�n�l�4q������.(�y��%l�3og���ro�Wj�;Su'�$&x�qo}��{��	^~�}f_�J7S*ՐBOV9�$���<�V��b�*G�R� ��N6���Y%���]�8�+�|rv&����R�ܬ�����_d�Rz��}8�S��p���B �դdYQ}���Ӳ�P��x�;<W�� � �=죣m�)]� �	}U���j�����p��ؠ],Ƞ��ҟ
e����I�*wS2r�YG�9hJ�ض���l�۲�V���NJ۱P~��"ݔ���%��x3��?�0%?G�
��\w%�9����5뗢1c9��c	w�[���X���׬,�^Jh��5�?,�@�!�}/	!w@�����E���{0�aR!��cܓ�F~x�I��Y"�3ʼ��G��L�R��Z��9swp|��d��%h���H�+�$l%�+�.��*�p�^�=��u�da�D���� �P�!��pwx_�f-KF�>
 �`�
)�� �@�,�T��8#����$m�.Vʏ������� i�r��&t�V�~��҇��n�=1��U�4<�i�~|"��S�3���0 Z>��?ʔ��C��=�HYS���_�X�C⌧�R���6JF�@��x7�o���-_=�Q\1��0a�m����(~U�(8>��%��Mi7M�v=���}pr�����&�[-��5��S��o��-�����Hr)��i�6�^�uX�xa�Do��S������\�Mѱ���P�+�
�I�^�^�GiK�
d|�㟭�Zq��x�|���o�9��HKE��]�~u�F��Ntd�z�s���?�����ҵr ����Y4���]�6�꫼�9(SҎ;���џ�M����P{a��^9,�]��&��]����m�T��������J���!�����<t��ڠ�d�O�l{'�HD������O���2�Z@D�	lb4BX�8�E%{��H`��6�K�<�y�c'�c�{󆇝_i��S���TaZ��6�v[8��6�yg���㠺X��aV��#ZF�SZgX)O�@��ό��Uz�s�̝|{]�x���/jn��t;���=��-WX�����_N1sN�l�Z���I/-Q܆����>�x_?�L���l�`���������$I����zѿ(1���[�6�7��C��W��5j����w��(��95�c��wx5x�c����:��� f�y�V����:��+b�-�����VH�����Û�u�  �/�5��#p"�L^0��*>�/	�8��v�P��r���'s����V���|��`$��P���D�w�:�@W�P=̳�� AG�����n�����Ta�eC��M���|"f����1�TzST�`a�B�|���Hj�^&�# �k/�-y.��DD��!")�ߑu�H�+�����?qL%�l���~"����n��}���s
]����Q���Ȣ��I����w�h�x?&��޿E�f���+;/��N�8����N:�@��Cr��WT�^�y�/� �O��Z6}��$�g� h(�s��d!��xW�B��hBXE�`���Y(�r.�dȘ��h`����\�w�!�M7���Y�߱�?�N뾝
zX�2]N��H���Bv½v���1����A�,�[1Qñ"Ӊ�`=!�*����M48$V\���7��|�I�;%թ"FOu6�$�㻩}��X:�T�C��:�=�}6�8�e-~����g>�M �l���X�"���0Nyn�MK���E�T��;#o���f��4Z��0SlE!�O䐓�aj�b�x����u:f��e���{P��{���wz���7���I��� 3�q6U�T}���H�"�'x ^y��Ik� g�l6B��PWk�3	<Y�`H��tBΎ�!�q}��SY��r�L]i��%V'~��
�N�.|>eּ�>�O�W��C���0��-�0�K61�͝X�w��%C��*��I���c���eLM/A�|we�2�H�@*�-;�LŦ�+VͬCW�[�5�U�f���[N���\W�Y��@���ɲ���Z��[�� �uVw��z���m�1�����#	�it��ٴkm���`����6*<��4X@U�����Γ�<�Ӎ$�0�X�w���~�LlG$�W���',�����1�06�y��rɵ��Q��Y�֬oܳ�s EVָ|,MF����-�%7�=K�ro�:=c ��ᆷ�����fG�����.���g�e����d=|RJ]�A璅��nLP�7m��<�?,��Sc�z\m��I|�
�Na/)�F��6D��I�&��՟#f��D��5�/���V:LO,kJo�d�d.��0�k���5T�|8��K��L��=�)��{׉�� �#_s�EA�i��0�<E^��J�~���$C@V���\S {�q�ޛ29�\����H:֖��a��p`�`X�P-���BE9�'�H)�5-��$jL�o,y0�u={�N������H��{F���ffqs���F��!��[��}r�p��[w�Bx�a{W���=�Q��f�� Q��$�rLT�;�m	Ô����V�D��LA�H�(��$8:Xz�+̄[o,>!
d?��!��?�1%�k�ye���+1��Fѝ1ҳ���w�I�fW�*���l4NE�|QL����#�;E#6׶!Z���=:��f'���T���+�j	0-�y���o�b�P�Qv��h�bk̽�87���^�.��x J��%D{q���_o��c�r�3m@�q�=.���T�0�����1�D���腗p�V}�V2�c+�����۠ (����������ش	���;<"pFI ��f��V�Z��8���s�T(��T��:؜V6���S�E6PH���mߟ B,�R_�QUɽ���Աg�?ӓ����,+8����[DlQs�.v��o� �᝔p�ֺP �l���	}f��9�h���-���������u�R&�p��|�jy>�)_���OPHV��$94��?�D�A����;�GƲ�Ň�3�~�a~(�}��N"gOA�"��V�H�H��j��+�*�*��̃Q�E�eǨ�{��.��%ʱ	�Cq}�+�;̚'W����Ro�NK�#([Z�)5j�UA���eD���Q{�u�ő�s��I~7L�D%�{�r���(曛���H$���qڪB�Kδ��f�Dz��v��'!�\�E�R��P���j�T��\�ȴ2	e�	�U���`�:�$�4��*CS>�G�`�J#�Ōi���I�$��G����2�V��]�%�SO˧ ?�49��(Oo�6I���lw����U��|y�3�;$܌���{KӾj8F�eD�.�MD9��f��.����):q��,3d'o�<�9V��\+��ĺx,���Zb����<�nă1A�j�"t�n�#��t
G�O�B7@`1r��.ˉ��}.�2b��i��n)W��0%#&?��j@�GG���'#��߸���te��V�U���lry^WѯV��s����u�Σ ���I�Ԭ�k�,�Cc����}e�\ƽ�е�����;�H�1@DcWsa7�.�,�*�H�喬t��c^�%Xh��z�S�n��u�Y�����́�����=4E��G�!n�&H�zŀ���{�O{��z�����	���Z���0(B�~sv�ˈђN�ѣ��f��n���Eʌ��Ӯu�I��4�V��o�_�Z� �$5�T�������������_.1p+���Mx�7/L�*RW�&@!��:¥>uv@,6G�O�)��=���������p���hg'�D�p�P�����2w��Ri{R� �÷��	jp��F)���:
r,>$KtiDZ?n�ɪ �(tY����q�n4G6�v��
C������.�#�v�ϫD.Ψ��{�����Xs�l�yL�V����t��W�����wmm'n��C��V�?����$�p�}^�%�����UE�ہ�r��!�����85���HX�-Q�[5$9
��(E	̪��t�ԬU޻_"�U(�K�N���M�YU ,e����M�i�L���-z�A�(�A���8cZ�9X�%�N45�1[�K���Oݣ��d���ne��`O�������
h�H{���<(L���-�n���	��5����^�9�]<+W��*�o�	T�_����؃�[�?Z���iO���a �f��:=�Tk-�v�&�r�Su�"�m�щ���ϣ�~>	ECt����8�Azԯ��rbT
�j��Xڢz�ӋŴ�������Ϫ����DN��W�TOM]{Snp��/��x \��P�k�
���b�]	Zy��^}��r�@���{���ᵷ\���p����8c�T$RJ��ZBg��Ct^�Dn�\Aj��=�e�U|k2 ��T453./ֵ?�{������
,%C5���K6
����{}X�<�(�����b�uJ�D8&8���v���)���k9�UF:.��W�̭@/9"�e�/ٕ?2�HW-���a�ʽ���9�6E:m8R���s']BJ��،� ��6]蚚��R�+���"��'��;v�0�N���5%�*���&��A������z?�Ȍ�5���}��%��Rx�5��kz��6Q�ݼk���O>1jKspl��%%�C�����nZ�n�9���S���3��z���X�2ֲz.OE��d�]$��C����vM�T��:��A�~�q8��+���N��H�oZ��[�H{�vz�畜�%���ܯ�|ήO�p��
�'��C�
�����:WCwZ[��N��/�TÀ�[;4?�)�a�k��ų
���j��>�j���F�۟=ӟ�W�������_���z���jm�it�f/	 �H0S��E�Qӯ�1���f&ҋ!� 6$�u�������R�h.�]�Uf���UnYdY�J-�w,Nj�`�[�
=C����)�7����u;�ON�E}Ä���.�K�_!w{�<Ԁ��o�#H_��	��0��j9�X��,���q�:Ļ��O���0'����1�@+��$�mZ���vugw0��Z��d�=!i2���AL��2���.I]��Fp�u�@e�o9�hG�Y-��O��!��� ���`�:���G��.�Apv��x�Ps��3\����#�``��&�p���w�
����t>8�OwB�89�K�Mmt�l>�f��"�����'a�~���3<����Wy���+Q��k(���h�g��^��iZp�A�P�%��K0����`��2��Ĺ]*�փ�}��^�+k>wR�0V�8
/�]Κ��u�r�L��:� �e쳹�F�ԃ�G���t�F�T��Ơ�1�9��cCZr���S��')����gJ���E�+�lYI�L�v! *xK"��;\�S� ���k����;-;j3�Zx�UQ��UD뉄�A���L�߼�����ZԪ��ޛh�-�w�@��DX�o���uߢ�����u��H��B� ���ʠϟ>�j��u�[a&w�Ȧ+s[]�U�͕��i���I���^�[s���G>b'��*�y;g<=��ܑ�J��&�#|������ٲk�pO��A34\�%9�^Z@]Ɗ,a� 1���=�Ćp�_�bY�=Uk'�Zğaiŷ�UAɔX�����n0��]���91�1"�e؃��<�t02>	s]�8�o�t���[:�{q��cip�9�!d@^,*�����=��eǣ�����XND�ޓ$�¬����2���[�"c5ʖ���M��!�1-0Y}b�V5;#sGߍ�>�����T��σj�2��]�Հi��k�`�}�)!)߼Mu �<	�m���c��3kng�j.#Ia��	p�,/(�K�,=_�G��{��� bj$�oK�"���koY�C��3�)//S�S6�8��%�>L�f@�Ǻ��ٜ�7z�Y1!%nU��*���E ��Wz�p\�O*�	��ʜ6e&}�f�Д��؂ "��g�φ�j.�4��K�r�y���<�"�D�/�<*�F�2��ͰG����/����)�
�A��z�.�t���6�)�e���Gf��粁r�Vla�;M��8��nk;ܙY;�Vtg�Dh,�C^����=�B��%q-D��z������P���~���Qw���6��0,5\d��G/a��\1L6�-����d�b�\���m^�ejZn�w*���-<�{��گ��<�G1�s��uZ�I�(>��RҮT����YoK5�K�f{q5���\���Bq�L�F�[w�N7��Uӕ��a��gu�o�,�7����츉1UV�0��;�K��f��V(�</�����y֗v�������N�y���|=:�+8y21�A'.@�O��U�P΅���]{�G6�����fG	��~>��:Ŵﮫf�5hX���S����&ܼ�>/!�V�*:�H�|ځ��l��3J�3�e)= nF���S�xF�4�÷��D�h�򴓀����v�d�R��P���i.��W@��Ǯ��ބ1��nR�E'��A:���+�Y�1��6��_��\�����w/; ���l�-Sk��7���spl���L�������L����Յ��]aA���A	ΨD�m^G���(Z���>O�,�\���B&,
j*�JP:����G�#����ك[}�#���D���@�g��5�I������B�.��譶O�h��T�kǃ��v���x��Զ�zS˛#zNm?3�f?���@�W��Z�^L�8
���M�C$?n�W�m=3��yn�P�M�+�
Tu����:R��OcZ���Y�Z�%8��;�ّ�8�;.z$�� ��������Vs7��цt��v��p�Ȫ��O�i����ы�N�I��\ӯI^����ȍ�2�'ߋ ��ћR��w�[H��)������o�0
�o�:-Ǉ��N���c���l�#�F����� P����,���G����xU����w��2��չ��d�>|R�
���6��f�vƄ���Iճ���Լp���z�9�r�i����q������z�}�"����ǵ����4'o�S����EҶ����	����=��_��lK���E���A���h�ud,Z�fT#�\ 3����Kyr���.�L,<��ccd����~3�����R�0�u� %6�R8�]����ɕ�Z#W�J+.��X$�Nx�&;��Ć��(! �V�-�:�C�DD�@<�.Y� �
k�A��ٮM�Q���|_�ی��_�&��3J� �@�0E��ݮuA@J�����j��{�?��@���m	߳W/%xO��A�XPy�H�a��Ǻ��njb�8-��M��9�a;^K���@P6�����b��/�3��c�f�F!�P���ʸ��}T�ώ�^��Y��h�I���Eo���YH��~�	&m�ݏd��M�g	7٦�� �P�λ:��!�\�~b�P�@�=ʁA��~va���P��K�&x��<�����g�*�b$:n�~i������	󺍀�x7���/i�e�s�Q7/֫�6pYmN�:��i��ڔl�Hp�	�}���R/]!Jߪ��[���[�d[N�Ll�#�����L���h����ʏCy�f�� qj��-}\l��p9i-�8W��Y��"���{�D��d"�_�7�(X��F�:��'�<F�*]Y��������jCl����P���d�U|�Z@�bCԱ�;�ڙX^��Λ���!�I��z��'������ ?4���D��z��7�sc�Y�}�	�O�i;��K8���o�Q)�s�S{�lC$5��T�I��w��o3c��4̭����|a���Eo��r0���ó8�Y
 �+
�'�|����~6��
�WoѲF}KF���WF_Ʀ�S�gh��
?t�a����oX;����-���<V�>%UT�h��J;%���X��K�Z�؃����.'��Wx�����j$�����<h1�W�#�S�C�=���܋��A\�M�E��I+\��nrkY�e�5 b�'\��k,�+zo&݅���5�,�E�.����uvē�����<���.��QI�1�iԻ:�l[�fՍ��|�z��cSV�G��F�x	��!%���f�a�����Ys���+�� #�ɓ�F�g�`sl{���\�a4�Wmx@��ۖ��f"G��@�E�_o�dA��}�P�L��c�2o����b8C�;+0�pm��&��~���~�Ì�H5ҀM�[�+'��1qpʤ��L�P�E?�^�L��hy��Ѓ�ʝ��+@e��ds9���������1��AJ�l[~G�����xnkP)�h���K��XQH��Ab��̆6 ��
�p���;�?��8F�AA\�<~�Ĥ͏�烕ĽKǷ�P��З�t�`L��N0�t���I���p(�%��x�ffE�4�!������p$�)$VxBd���>P'��J����h�>�'i�*�g�81
��3s�N�D.�B����tT�{FB*ͯ����������ʻ�km0�"��e�z�|�$�
�M0�ݸ}h�e\e3~�|H�ȩ�A��Ἱ�I=p[�/3��q	�Q��,��yF��nCnBX�@|R,�a��3[�ټ�3)�`YuԹ���Tnn��9E�u*��;��˖����� K��lꐮ4[�ԟӻv��*�t�v��ܧ���9�2��k2FJ���t�+�)+�ۘw��I�_�>���ۀ"�0�} ԙ�0.SDV�["��v�K%��_�5�O���AW<���ŷ��+�0-�+�o��C����?�T�nU��a��}y@�\R�ĭ7��SN�,�8y�A�[c���Îx�� �IF�_Ǡ;%�뫆�:�R�᜻���P�Jxb�Ј"�k�C	��,��Z�Qg��k��٪*USc��G*s	���k �0)�3/�v�*N6C�����]99:"@u�h���P�M$���X�d�8t��-�|�d)%���@=?6Gk���3��:N=Q�el�S֭A=x]`�h�K|�K�ds�D��s�a�+^����W�+��d5S/xzܖ��Yc�ie�z��̚�
��,5���"N0�����XVf=fo�ئ3i�1[� �?K��]�\Yz����h��Q��/���\����c �5�[u<�*~H�.<&��6L�Rt��oG ����K�/�2a�x��є��(�TH�˱+.(��榕�s�*6f�ͮc��-%�y'�*�<Y�Co<O�t��Cص@T�	�\̚�o�ëD�a��[#��s�dh�r(�w�AS��db�`�rS��&�w($�Ee������W�=.$�UU���y(���	��Uu��&��<�`Y5���*�J�fv����޹�Q�@@~꫋�2�!uy��%SB`�t�G���� �����m��"�{I��h0�i��<�]q���T?E|3>�i[t62���x�S�4RM�5� !�f�I���3�5�ܝ\ϊ�l�=�%GJ��B6���Z��R����}X��(�s9�zɻ@|��_�����F9������Vh��s"�d�2�b$��ò>Я����B�g_%�޷�[e���<��%�M|��0����y�ғib���v�|&:�!��CP�D�0W�͵����l��a^�.�2z?CѴB�\�d�����L��8�����Ї�
���T��ծf5�fx#y|��t��p�X���Q������{����%��+�[OѭiKb�G)Y�< �S�x���(v7��{�?ճ�U��⽞s=�O;��0^��}�NLf���v��OS��_�I�U5�yR]�(g��%p&u.��h3�(��ѳE��$)._�Cs���c�[�CY�޼��d�{#�gX��a;
97%��:�����=-̭��#Gd���]B�NUL���Y��2i���B�N5�#R�a�ހX?�7�3���#�57tE����G�œ!���Z"����$���`��1J��<�X�!P��6��3F����8�S�*@T/�ұ�]3�:q'j�<�W(�S�m��y�S�VF&䦒���6h�Ǯ(	��i]^�!g$S�Ѥ����p%h��ړ�u湭��K�^�*:x�p<.zy��9�X���o�+��Ukp����?ߍm�g{am�yJ����NP�?��C�[9kSC��9�$P�rX���ӷ�U6>�Fo{M/����}f�s2��wj���n��v� '�Y��j#~��I����SW�(�P���e���k0x�>�)Cc�٘�M�4�������jF�6V�|ɐ��I-ԅ�mP�}��އ!�պ���������&o�d��KB)����D��i^��#�7V���Ղ�`1v�����8;�Z����@��6��ר?�l��
2���ڥTpg��+<������1�^����L�5X�.�lw�N��~h')�U��[;���=bk����e�6q��Y�
��]2ï�j#8��TRY?����L��=F+;�=(��U�N�%e��3������sW=¿`6���l,�P?�J�v��!��Jz��J/%#��+��Ů��% 2}=�bL:�>�kF�r5=�̂ Z�9vǧ,������$�X���}�u�O�&r,	R���5���<�ݸ�����YY�4�
i+���,����l��`m2;3zifE����U��AďT��~�=1���&a��(k���B(��W��a��A���J��F[8��Q��z꫁H�.�b��@��/n�+4��Vk]�=`����	>)H<M�a6�����O�y�<"�R��}z��4��j�H|]Z4���E�l�=YE�d�����+8�J�@w"�O����\ �E��m 	��f�8���l�btT�zF�ᨒ-�h�M� i��|#y�@DB���ާsU�+89-*�۫��z��G�z�?T� ��r˕+W(F�x]��z��@��
ַZTz��
/+*���SH����k��ɠ��ٝ�S��j�a"g�I�j2m��F�J�,�뎘���U[��x$�uA��c~ !wko�!�\���i���ߑ����o���6
45�h�}���<��!p����������菺
�P+H��pej��b������y�z��N�?g� @wF�hu.�����}��V9|�Mu8�����s����Z����V"���%�q����	5T�4D�)L���n�<wu��̅�HxQqR�uA�&FN�	ֿd%�	:�����g�\���`�$����4Qo �n�u�d��e��k"��ƄgEѠ�T��[�2��C/���Z��9U�TO���Ԗw��ug��l9u����~�C�ϜJ,b�>5G�l�3���qL����\�`S��B�S�o��d�gM�Z�7�E���8|ްSR)~���N׿�v��W�*������_�wi�����y��^[��L-5�u�ڍ�9�I!���V�j�=���w;�E�Ri��]l�����a��>"\8;._Y���v6��Ƭ��Ix��s`uK:e����rs����$ת:��!Rރ1�[���	3�N�ͬo�HT�Rѯ	���^R����}�F�4N4fȟ�Ra� �NX$K�Ex����jS���P|b���hХ?/ �+VF�Ф�yCMWj:���̙�x���~�������N�}E��1v�ړE*
���/[<����F��?3�:��h�I���<���=QP �9�J�VUĸ6�⠭����Y���0���Kզn�"u.�>6[mr[Nտ���.�E��]�U�P�4`�鸏���Sڷ�6�*���Pl���"�.q<5��8Z;��I����BCp�F�ך8�{c��	�øv�6���{q�H��J��{_j��w�ϓ�W	�)҇�Ɗ���!o]JԽ���w���YbD�u������Yx�c
-_������K����<�jC��uZ�f���O7���Ƈ��0����3�^2C�;g�A٠�S��2n��c::Fq&{��T�|�5HoJ-��a)������޽6��t�g���鸰-	3���@�s�I�5^8=�q��)���ۜ��x�v�%B��u3P���M�6���_=�d�-+lr�������-9�_f4���:"��er���S�K�0	9����9�Ģ�8�u(�,2��C�7��8�����W��'�L���g���w���`�-*Y�cU�;�QUѫM���2�I+.����݈�u�� g�k��Fܼ�F��73�����X�s��y�͐�Yߖ}�g0�X�$�=<�J�S!�5�uL8���B'�E��<� ���*	eC�=��I~W!�7�� �W�[bZ�w�Z�tqz�Wpz�����)9��`#����W.��Tcj�(����������=z��W��8����2�����&s��g  ~�\a\��'�7i�Ὃ6	����һ~JI�/�$v5��\~D�ͼq�_CvT�t!�$Q^Q������)%no��L|Ҽ�ͥꩾ:3w�F�V�˹�_4��.<�z'!�cϘ��ĺ�~+0�����A�e�^�֔bb�}�"���j�[��QF�v�8'����k8�F�xB����nO��U��։l�E��)fE�3��$�Z�p�r���Z�_R���7_nB��.�Ԥ*��9�����n֔�t0����\P��9k�o�&��/M���>~���d��;M*y��-�/Ah���b����	mI��B\�J~4�����`�R�M�o��}�R��в�?���M�+��L�fX�۝ ��$G;8iG�/�&y��!F���G�"���#abʄ�`�����/�%vƴ�~A�� 2H�梒�k�+|Ĵ��$=o��	�!�>����?�����c������Gna!� "Ge�F�!�'����h$�=V:���xiP��5�mg{������CD�,��F�2i8�?�.�^��(�r X�'�^��F]���+LF7O�6�D	��G�2�84��@���^��Or=�h0*y�z_;����ߊ,��a�&�?�.�]X�Nψ󳛓ƶl�x��7��TO�<B�`�w�5/�1�GF�y�S�t�5ǋ!��X��ǇTqmC`Sy������ӝe�8Z�o������V3at�9�^��&�"^HEy�J�%k�I�r���[N ��f� ;�/ݜl�$�j�%�_�N=b�U�-B2Uޚ%�)��=��..����p�i�+�P2}S?݋	Z?���8�d�R/'����nlق��1ϼ���Dڌu������ق�����J����_Ҙɫ��Jb�V�-pv�Yx.Q���ucf��D��#��N�)�Ŗd}h�f��=K�@&_n�xىm��G̉+;{V���=�Y��4Pr�Q��m8��5�7���(���}w�*	����
wpL� �d\ }>�ZR@�`��A�ҵQI����K�t"F:Rl<��K�x�lE��.��7N�nC.hs�N��4����/�Z����s�R��t}4�y�߽��I= +ޓ/'���u�}:����p��n�	� 1`oz���	a�7 �D����3���'�;��#�W���쇁u)��n���m�:����B�.q�N���*$�C���3bbfX���v���D2�0t%Dh���Wj@M�X�!����yw2c�m�|�Nz�(<h���>5�z�]�'r�(�<�����NTj}��*�¤��f�^|3�d�N"T~�r<2���3"���/�# �1�2q�*�v,?(HnM�i^Q����d.W,�9g���Y���*�P[n�Z����}��Jz�UA�����[P��0c��K�Yhs�7���M���T�������K>�ƐrXF6~ҽ��RJ�>��G �Y��<:��U�k�H��\˥���33���ׅЫ5	��Z���NL���i�P�-}=;T=���ه�20�Q�!�x� $�Py{��M�B��>� ����I%�~��z�m� ���5�e��g�nM�f�}"��dF�3S������5�_�U�4�Fg�,rP�O�giڱ������bڇg��pKF��Q��%�����|�в,P�(�ɋ]� ��Q�v�~�$���?~�ɘEU8U�{�x�>;4�od��e����U$��,aB�s�C�T�����H|~EK�U�G���߼��1T�6�:���܏	$�4i>���YX\:��V{N�Np�1��Fw��I���3��-! 4^�d6����e�Uar��1:T�>�9g�����{=����q>��f͆eb$�'�����^AO��d��t������'5l����NsN����?�j�1)�ԑ�3v+�����6� 5ͻ�s���+x���K���m�ء,
��Um�޲�͐�j9(Q�[ �l�*,`N�|�H�|aAtZH��ÞZ�vu�y�����@����{j؋���P[:�*��.	]2N�Sz�Fi
=n�˶Jm�/��*�=¨�;d�cΣ�dy]V�����7!l:Wz���\��n���:�eCpQF�1�a��U&�nR<��=V[�o<;�j�w��g̹ke�`��0i*���<�f�����29� wL��y��$,�SH�����LN�8Yp���3��Ѻ9?�;8���
����qq�9+ɨ���ˡ�P�ܜ@el��|�ޏ�tL�+o�:��z_�0��2�f1NU�~FQn���u��Q��M���f恷����7'?�M�ǽ␈�ֈ]��
cJ&��:M����+���>�`�vE N��2��Iuw9���;�ʮ�n���!�TQ�T�!<�J&͜��cS�+9��!��?h��J�W�����꬚��6�j���}ct]Y��\���~���+4�u^�2A⋰c��M�brF��_M��]���94���(ʰ"Y��4��Ԍ�0#�z�dEڒ���,��UvA-���%�2��[��l<��� ��	~��x��5q���z67�0|^M�Ѓy�/�e�·��T�|
��<^Y���x⎳ �B�����`��>�n�^�O���U�I�����i9�.��z�FB�7'������n��ϲX*�I��>A1�]��sZ�ci��S=7)l�y�{���Xo��`��Xy��!냩:r������z<�q��Be?�_�� j�3U5�i�3ڢ
�+#h\��R<7����s���G��=`������^�RN��՛cJ�z�Ly<�]�n�:7��ҩ�l^m�y�h!�=�alB#>��s���I����<|��5������8�b�9z����,L^�LD"��K.�:/����λK�֛�l���_�.�g�T������P�֌�:`����_A�b�T������V�w���6����c�L�ع)	;���F��@�ӕ�(0�:��d����v�*�G�.|CǱ�u����s��2~л�\T�gw��8�UJ�������'tm'�Ơ8��1��I��'�P����H�AI)*��8ʱ���ހ�2�>�+�:��B��H�;��6A��;<ؕ�F�`lId�/ն0�kOwC�����!5���J,��5O���P��T]���L2�)�����X���	�@�MV�|�</
K�n��(oL�=︙�p
�y1A�h����dܳ��+ʜ�`P!گ���S_Z�r���@�j2�X�sМ-����?-	s��`uvVYv�@�;s�O�(�B)ڀq�ő���mM���")�i���Pb	w�G�?�B�3Jg[���F���"]�s^`ܮ0[�s���§dʙ���aû�����r�_K��z�}��Y�x���%85�x#Y�b�V�F^$#s��B.�ȨH.�W����Gj��+,�+̍��t�n����y�'!�J��St�b���O/�o�>$�W��ue�D�<^�1�N����N��K���wi��)��T���C"�b������ ��][��� ��%�J>@��
B�_�Ll��<�ؘr�ȳIݡ���':��;>aj�aeD�D��D�\���ST6�TM)��m���Չ�����=w	�����w%����#�b�����t�,
ŗu�&�Pzi&�I�ɬ�Q���[J��K8Ƶ߮Ō�����[��k 2���qB>�W�4*���4�R�"��%NX�,�F���w
�0�
��|k�s�Vv�&H
D��G��g�h�,�!s�}30��ª�e��-��E�Ҹ������&D�&��V|K�d�o�ԧQ�,�M�:O/�+M5��ǦČ��y@�eq�ڊE藃����*ТH���]+������� �jǎ��SPn��0��Sg~����/��u��*@�����/�'J����e���?����IO�`;5���sǘj�-����޿qN���"�!���\�~=�u�}�������#�U��}3;c��g�z��*���>������?uA�*V���¨v��3��7o���%k�Bm"Ay�o����-6\b�C�Oӟm
Ζ���4�Ã�A���#tl=Q4J�66��._�d� ��CO��n�5�����f�>'�VW���B&�)���.�00�K|�_O�A�a��^h�Uhr��(�TJ��A1�@ܮ��r��ޚ))P�*�����X:i���u:@]��b߷i��vm��/�(���1��c5�<��$�ݫ4�.�*]�:AR?���	i�u���t���œ�ݐn���F���QKj��J�B�-��e�wd#�a?��3j��B�6��5x����z�6�~�R��lmu�����\���s ;�NB��VIĭ�Vd?m&^�zNz��l�P�� �X�|�M��Dr��^)A-��i����>�} B/��@.�ErZ#���-�q��FjO�/h@�bzc�''Kӟ�,Ch�FWE`�᱓��!2#��F0u4&���T+�Uh���H<2_Wˏ`����S�\���^!�ZK�E�r��N�}��IA{\_t��)rd�s
o��_����j���Tb�N><��,��'!F^�Q�RDmv�X$����m�WY��X��1 |l��u�桚�j��ι��r�#��J��P���:�vWun��C�4�]��Ǝ��GC�a�_FU�Z5kc�������n��Z?��Kl�����(]��Qu��V�GV��[m��U\ε?�LCz�O�,�5��yq�B��*���`U����/S�Hz��>X��{�r_ߺŝxw|{M�v�}6nڧxwZ�Cy(*y��쯌���T�ߣݔk�0K���p���h���+⩍C`E�0>Zr[)P�����x }w����	��C/�EØ�����]2l#���v�����R��Mѫ6�����k��9-�Zjȹ��l�B�%��(<���r���\ �y���X�OT��<��������'�G�K�o�:��1�4
 E�3�s��s#������o���P��^%��}b�EA�ߜ�wp�8{H>�[��:c@H�Ԕ���4]��9w��UȂ᥸>��Σ��t6`��?w��Z7u㨿PRm'nN�	|\����_��a:t�(�G<b����e�����	�� ���B	�����ٹ��T���q��;l�~R]|����<o����늙wE���u�0f�:��"4rظ�&�yK�+�*�n���y E�'�N�04�|�l�_i�U�ص���rP��5�B���4��_?@����د� Lp���y쑾��?���  F���4�L�����]l����TI�I���a�][v��E�&�CMǘ��p��$�\p�����է�(4�#�%�'���R�٘�9�҇cn9��Y�!0e0�ڨg:�\��6$�Y�����d�t]5L�	\a�s����Iy�U�o4�������EutrK���̵��Ñ�K�c3IR�_ؠ�i���"�ߣ�D�����]dK8�zm��2)f9'T���ǁ$��9�����c[�jPn��5��E���u�m�C�o-	��9��ѿ�c��_���?j 6`V��j�x|�g���l�@|K��˚!G$�_ƒ�G*/DL.O�2�p�P�&�`��!u��F���wiע���5��:Q~�zT���z�fM愪X]���>]UO��iYN|��tEm�]�E8�>&Rď�mY ����ya���i�QV-&��	�C���w_��P^ݨ�K:�׾g������0<MǏ��2��/��9�����u�գ�Q�k4n��?[���6k�b �ԍ��Ƞ �>p�tY ]�6�Vc;�1צힷ�oo��q�Z�Imz�4��d��>��T��Fh����y=�@l��SO��Mޯ�,�V��D@��:�Ɨ��.��*}
ZAr���c��d4(�j�Nz�Yһ��C*O�E�w�t�2��O���P���j�6?�VP�����X�T�m� ���'�u�'Ps���Z��� p���5ц���Gg�p�x��/��Ky�����,�a��H�h�������t���u7ڹ��k��"�l?����,��$A��"J���9#���Q�ݟ�(��]��
�Iᯏ���z_
��#T��'����(��:@lAVHs��H#{���H�)��6�k�1���ߟm��9"��N��"['^a?�G�-k���0�v�T����F�4r�"6%ޕ���6o�]K.h{���ڤ� �C$�ys ��ŉ��%�m��A1�٠�
�|�)�d�,?���6�q5���pp�I�h�C}9(�J����j؜�ʍ�3���a���e��zŭ�T�R�`������V�NP�a BKH/ޔ^6J=���p�lD����[��������`���)ki3b�h6��%��Mucl}�'Nt���`��uX�G��m>;��\>�������_�	���<�O�i*(��R��-I�V͸%��Ib��0�P�k�a����x��2(�nۈ���=tT����[�3����i2ڂ���AK���'
��$���V�hGJ��^<�gg��}7�Z�v�I��E�N�*+�N�IT�L����0?P�}��ˉ�ncWOu��-�I3K+��ƴ/
n:7��d��~j�{��0�W�W�y��Kn��9��k��(��]���ؠ�}�Z�i~��k1g���^�jV�ZҁW�*�f�#���nVz��'�Z��`晵t�6^��ZI��1QK�6o�? £H��]�����F��YL�b��R�Ā���[��V��Ǆ�����TB����\�+����mCt�D���ߨ�3+��w��"�;=��N�)Mx�0 O�����d���7I>��:e�`]ixw	޻~;g	��'m|]o�a�,�aDMG��d��Ɏ�YI`%���(��lճ������a�<��;�m������`]��h��N`N��>���
�{�d���@��l@`���(ժ�Þ�fL@w��h��U����@2�ԗ�^��9������"��>��H��w�u�$�OL�M+�0�i7#L
�QN�i:�Q �9��-ՔF Bڈ��%�ߕ,Ϣś6�<i���#u�����$����]�y�`ח&5��3&]��v��=<[���UY��g嫿�gJ��~�?���"I$V����M�"�t��I�9�a'r�(7��$��?�W}�1"��ԩ�F~�G^��G��j�S@�*ߜ������KIM��80���< H8(�-�_����/���}�sع�}o�F���!3_��w�7H�(�}E.��PˣC�~���Ml܆�h����!*i(��"4�sr$ǔ�*x����v���]�a�l�th�#�%Ȓ�1�)����	��i6cN}@FX��\J��'8��D����i�a�G�u^����D���W���ʔ����DF���:R�؈S8��pC"dC�tu��/��QD��So3�5����R�-!���-E䞍؞�k�ph���:�������ו��g�{/����Q�����C#�qe��y�5.�S5��\G���8�in꠮,m?����x�#����& Q
�*�K.k2.�/z&��nC�+C�yM<<=�o����-I�oI��N�#����U��T��
���vzV/�+�C|��d��aAOF	���M��{��v��լ��g���aC���B�&TN:]go��+NN2��=`�D��w�H�.L�=jmK�u�:��+� �����D�0�'%�{8��b~��o��8:>{����!�jL �97��Iw�~> �ٵ�[�$�'sr�A���A*����<1�3��Shi1\��k�P[ik�m`ly`��&2
ĥ#�ǥe�q�� �X/�pag�<w����.Mw�vb��8���JB���.Fc(�<�E=��!P' �f�{��>���X�t$�+|K{�I-��fwy�+��G�F����C�`���q1���w��A��k�80yeI}\\KH��|n��Toyo��P�aIa���֛V.�^_ܘdTT!��֣���G���.��/uT���.�r��٘� |"z��˓_r����rW   ���n��E}��qt����`�ւ�P<�0Ƈx��v�ێ���r޴�� �
m�O�����Ӱ�Шն�t�;2 h?0D�Z��/_�7!ء]z��eU�<'k��Ad��࿙Op�B�%������� [������T�s�p=nՑo��!Y n�M����f"0��^��T�_ͷ�6y��t�w���c�й�@�75���).[T?�X���*��r6��#��1�¦�}��D����0�	���l���@̟/έ�H0S|Ʈ�@�ƒg�0MEs���J�6��1�&S����I;����v����U���,�չ$� �W�0[ �r���S�i��������@�ؿ[
+1���O��ߍda|Y:��X�w�ʇda��3َi�E	�+sp.�m2�l��۹���l	�֘t^d��>|Ęl.X\q������ �7�@����j���>����;o#�¯��Dk���i�y���6�k����jq܎��9#{?���P��ޚ�{�P���D��2o�	�i&qkw�r������-r���	���o�9��g����h��b�q��J&��|:N"����|<X�*5�Us�HkSc4��ٱ�`b�L`��ʯ�'Ui~?4�1����t�-3V����_a�Q��줐�o�8m$n�	�6p�^
*=�ۭ�\A�5d��O
T�7s�߄���
��t���	�:�����U���$�Q&c�����ݍ<|��!B�Ȯ<�p[�D�}Q �g];�Q���HK��sic�CN*�uD�MրG%j���~��y4J{�BU�U�j�S����H�r.�h���_=�Y�;�(�z�nl �!ܗ�d�N $�KrE�S.�=	z�Π+qWQ3���;7����(-I�AOR�.�K�4�/��> �.�����Dx��O�*x:����Ą�~L�	N�{o��{�A�Flq/잟M�����
~QFx�����~a��ZE̼+V����"Qҙ�Z2񁺢S�;�S�Q���LU��@1���c~׮2�/W���?��i��/<�-����r���o��3MM�H����Ff�穦�9� �D��8r�����I�W�P�����@�lpe���R�{��oX�F���5��2qiC-*�E�q�0f`�h�m�f�SR��)!�C/�K��Q��!ef���@����"��o%u:���>#���*��M���&X9s���@�=N��m�訇4���֣�o7U�/wk�eF��zi)G��I�@�p<ő���6@9��X�� �Y�bb�� l꣢-~����(rP!e~����gq�v\As8��9�+s�]������a�m=��pN	1'˰���N���\�k��ץ��pVDXn=���8�c�KE]����:�K�����#�q��&ʜ+��M2$��]/&� ��q��81��턲B
�'4�	q�F�L@�HV� ���W���g�3���Hj����Dc�X�k�~�&�xgLpO�&��]D��2�<q<W��tp�D�F�������|�Q���H�݋�J/�16�vR$��xAo[�u��=�FZ�[�9��p���y͡`i���*�D��G�z�&~����0�rz]��Ab]E�m�49�?f�E��W�ъ��Gb���nn[r����Qם;�m��D1ul�!����f*G��Tz�<��iE�H�u�:�P*����E�^�2a-��T
��)�Q�GE}(� ��]���p9�ua�@e���O�f��{���Ӻ>"[Ѧ����Fv�S�j�BYs�����ގt�]��㹺D'�@dzt�`��*��l�r�F;�����W�k}MdK�O�[����VH՝�2JM��h�j�k�ŊU%ҋ��M�EVg���rw�+z�`�l�o��8� Х�#�ϧ��4}��
%��b�*�&h�������|�N�� �����Pn��������~�
� �ͨ'4;Z'�_�B�=P
E���m[���VԛSRs��mq5b1N��:7J��j)�=?�ˣL���фC.����Y��? �B�d������ ��]4�O�dB��l8��O�x�v������=`�W;M櫳��#�ȉ���t+&��zQ-*�~���)���m�&�L��1&j��\Y���kVڱW��R^8x�q灐?��=������^��L>�0�ȶ8��KmA:R�׽�(�l�:�V3F�r�"N~���R�qi�~����(ზcyCB�>�[�7��vY�9k�Q���\G�K$���_�i19����'��N�f�ő?�h��U��w��H_Kc�����YZ�)n��f H���6��w�p�E[��G�SH����7	��8�̎5bK	Moc�q�^���Y;Rm} �_�q%Wv�Ah���L��,k�>Fm �䰧�1�+Ā���3���xu��R
�w�:{�Jg7�k�X��s��&/�r�KJ�G�"�!D)��(v�r��Z�_�q=�Dki��<?T>q���Kv����/|�,v%�v��e/��3�C�M��7�q�$��XK��ZX�����Ɯ�{W����k"%�f9}��Wx�ީ#P��.�lb$K��_�[�8��d�VC	J^��Q�H�[G��X�y�ϑ#����0p��Ձ,����/��,S!nG	)|�|<!���n�g�����6�0����jj�Z��u��^���>N�ο��@���$�t����%������A,���˸�i��#O��f��)�#�t䶩�unS�\�?[��k=)�)�d,S�	U�]��]��L�p))�n���3�j��%%��S+��D�%`i;G�Y�s
�@u��d�:;�c=�	�4����cӰ���
IK���!��[���a�|�*LS�ɬ��ￅY_�w�ۂ����z'B.'��2Sm��M��g��3�]��H�"�J��&x�0�mh�^:
S�=�.w]dHé���&UΒo��Aih�\5�]�"rf�
��j^�E�W\��a+V�P�2��Σ��o�F�'�qV 13x����v�"!��o�f���`�֙G ��Ӌc����	p���ԭ<��R�ŀ:�{����oO5�@�>ώ�(�*)���*w�e�C�W���,=XPTX��yM���'Q4�1��N&���!9@��Ζ�y�fL
L����+����8�7�"_��/��?j��
�?KB���?��`�^F�����D�7�a��)��Q.�d��ZIcC�ϋ�Es)c	�/0�r������$s،�ACI=�R�^�V'ܕ���� ���T���Z��GF���G�jx����^�{@�K�E�]��C��Q�ZE�#��;m�1�Q|1U��q�-�����3��,�����I��(���`�.��` �)�v�M~L�8OgX� �> �<�,/�lӤ�K�CfVuu�^�q��H��k&Im��X�W���)���o0(���N�o�+�/�Cv�q0�:��葚))�x�0�m��+�n�� ��r^�<���#�]/��j��;,�RKQ7۶�Y�K�	%����d�$D���w���u�4]T	0�l7�N�:��IF�K� ]��A��8����/P��i�Ȣ<�[*�/I��uęڹ�5!І�5t��Ѵ،��
,Y�'�4
hG��4d؊�� �J�ul>g"�DPN(,����i��K�.�g��_�ġ/[&W�Bz�jZGѲ9(���8��x���M�RB![��M��ś'�����v�;}d��Ij:f̕�B ��� �=�����i�'�G��0���n�d8O�	'����	8D,�GO��(�R(w����NI\��:۝�B��2�?0�?�7y5�UΎUT����Mp�q"��-E�ז��wA�oF<��[�}#
xN��/�xD�#icy����E�zOq�
�\}���n��,?�9��d�� ֎��������ѪP��>�(&�$#d\ ɨe��D�,n�0�Z��K7�ԩ������1��r����7�سp��9}"��:�e@k+)X��]
L�R�Gq��+�2�W�և��sh�B�،%i�s�f��TJ��ǄVV"�x�A��_���b�ڣ��I�>��Q�ߣ`��a�f��?=��M>��o=wk��6�?�Q�����<��R�.������:#O�����/��b���l��vv�a�����^3$�[c�B������&�{Ծ�>YA��jxag�@��%
�UK�0̵�y�5���(c_� ]\G6���!�1��ӳ��w�=��� Bg睱E�Փ>ok���R�;W��$���q�!���h�����N�N=�ƫ��"(_X��(�p�p��9=1����=g�[�u�f*=4��M���.G���A��=(;���/"I�_\/%�X��2�����,s�Ԑf��ؤ�W���ܛ(o�� �6��\u����5ҩ3���������I+�wk������R�=���"S��C7d�_�۔rD!ӂ�ٯd[���s���J��5�,�7�*'U�1Nh���<�A��{=��t���p�-��B5{������AB���m����e@��]I��*7����DϐZ�d�DW4	��lgA�]i�9Z��a4`l���ŧ��a-�	(�����C��r�*���"B�~�
8u�����[�җ:ɻԓ��F[��sf	��2�~����ല��kK�6�a���w���,y,�2�c]�{k3�0�����S#}���9��SeS{Vln��h�)D0Mp�q����Y��lB��|�y\�� �,�Z؃�i�:�4@��Z��W����('SD��?�Y��mX��c����g����
}�e�&	eW���g�榯)��oX���f9^rq��bHk(�b��.�{��4I�����lОa����]+˪)�D�辠�0���\^��J��SN�4T�(ݬ���y��:[��¸{�_��`�	Z�Нm�{O����z�_"�V�>�y*^֎H�bㆆ2�\��)(u�"��A�� 'XK-���|ns�j��ttK������#!`���+����ѳv���~��f��v ��������<i�SXz�/��Z=�PbD�a�	3=ӕ��R�
��x�~�B�x������яXYu�PL�P@�c	mo������^�_Ѕ�l����b�@G�����t�xdDHTi0?%��4�y�����s~8db�eY���tW�SY��:�.ѳ��鳐�~C�!�����a	��f�g�����mԍ��<�=����aT��c5���C����^��kOl�[Ɓ�w�_�2�����>���t����J��C��r4z���;�Q�H���aB��\!=Ho{_��d��|�oq�gn��A���W��*sk�N�^�r�}⷟#�.W���%�i5S�T�rh�hkcn%�A�Nf���v��Q�g��ǳ�K����g��-�����l3C;���ο�_<�>�R�(�9�1GY��^.�2N@35]�J���z�w��dtO(������|e�C ��r2t��Q�M�+�IA��tb�Eߝ�=�s���Q��L8WP}@9�)�o��p�j;?�U�XxY�\@;��!�ο��
�+՚"������x=6s��'.cXC*�oXs�����~�f��pq�u�s��ž(K!Az���ݼU�f��۶d�("�o�z�%���f�žҸ�P�6�E�Q���m��/*��"����[S��i���iK3d�?�s��g��=�_�]�'��eL<ۜNLӻyB���u��k�V��R�M0�dG��kO�&?��=.�e�B7O�bѮ�~�}`�C�C&/~M��o�������Ւ�Q8�EX�-R���0��K��=�v���jɧ8z�L
!)���kH�+;�"�N�."`�M�;��'���OᣜH���Ce6��i�q�~r\{�NxlWD��7
]�(�ۘ7,WB7���k;	Kۜ���@C�C��yT~K��I&���
X�IŘv ��N(?�	��0V�dݝg�J�+�#ٗ	�a�?��l���A�q��s�R]�ޏC��z���RmB2 �B�疁���8H v��`��;���j�f#��Ń���ES�n@2�� {4A��{%.
��4zlAkbX�u����ؓ���-�����\�*ß�R-٣�f8ڞ4`�(�-Y�uհF�UǗ~�UU�	���ư�GQ�ڍ;a���F�cp��8m|�&@�rS�-6�H�%�r�F��_~� 3�;c�u�+K3��d&\SG|�s���Cay�^�	v7!
�,������[�I`,-�Q�Z�>��qAO�1e�	-���-OӂO� ��"�)����'�Guõ�����M�2H�S*�$L��
�x����l�n�	��H���g�p@�� C�,���?��a��6Ǳ&�l��bN��1�O��H"I���r��)
H���W��L
'�CG��.���Z24yG���mf�Q`uD�L;�������j�8�J(�3�}�ח;�)�3Z���Ns_�|�s�v]�/f����tt}	(�c�����ɣ�R�W!N4�T��N���A\}+��GǗ�u���!�j��_�����fY�����!p�-á�Ξ����rЀ�����&|�AG�O�K�%���cg#�b�.��nh�kP��C%"Ǒ�]��`�n9|l�L�zo@%�MPx���m�A�Y"E��VfR�n�Ӷ����v�ʰ�nv".��Bj?x��A���/����*�s��{�+ �d'`G4�>�<�Q(@A(lY���8(��xs).�;���l�NX-|����e�w��c�~7���MwΑl�S���J;�����)� �{�� qW}�$S&�'��
����dJ_3�%�`Y�hM��$Id�NԸ+�J�	����O�4��ҙM�}�!��˹��+�F�*h:�i0���=%m?��2~��c�S�"kA�g]+�j^�������Q�wθ�( �yB�z��vp,qbD�d��V%�Y0�ay��&7�Trv�|�+i4!�w�Aq�"\�XJ!�N��P��}/yn�������Ao+��b\�'g�ĭ�H(�Xl����Yc��7W�;�$�b��Pz�����)} �:���U�t��U�I]oM���#ZQ:�0�K�Fhjg�X��:��w�c���;�-J��C?��e�vl���ىЃED�m��v�����L�$�ĢN�0�A�;Szm&����q������r��������i��(B�7���J�w,�8ԅG}�� v?�C�:!{�R9�0����,��)@ ��*�7܌xѮ=��W�bL|%b���M/�� �q�W��S��}cBj�ů��D��a��$�%�q3Ӝ�c��;�F�~��[�A���f�X�y++����m�t�c�a�Aqϯ%��sd��I�9�nR��x�A/���5�$�ѿ������+Q,m�({�n��5��2)�^�H�*�J:��4HBj�p�C���v��[����7 P�����X�g5.�`�mK0���Δu���\��	�F�b	v:�v���2�$�{х�l�Ў������(r�\
/V�R!�7�����P\�*�âԀv}+��CM+i��G��/n�
Kal3!@�"��v�[|R���P^2�G�W�p��Dp�HT��>j��!�8{\u�͍R��#p.7�I Q��~;CUZIz���x�`V�gyN�>TN�=�k�WF�w ��z�j��<�����E׿#2�͋Ǆճ�~N����nvF1����Ӹ�*�ojh��+El(��
�c� �mQ�"���O�����ZJ�mv�Z��H�b:�j����χ����N"�c���&OCa�
��wZ�-�5<�ks�s�A���YЉ�eZ�.L�����i����/?���ۙ�
m~�����|{����M]�,r�Y^��~"9忷N��W� �*����[��F��e����<ӱ;wI���jTuG	��]�u�̡˭�40�Ώr:V��~+�-��oj��a3\�)��A�9���U ��}���F���4��!�7���(֊d�0��7�=� YV�h�Q-��
'=!��&u �(#�5Y1�Ӿ���b�S��*�+wcE�Q�&/(�,�iu���Um݌��7���<a.(����3��^�h��'�®�,�.��}�_��gI��Yz���!��s����!��Kk��H�Q�⛷)�2nBC�-���nm}�ʐц���X8��άZ��ap�\�AF����!����b8-�P���������ecn@;KX�O��;�W�z�~f�i��Y맆?�4�8� �R��YG�O٢�/�V�5Ρ��D� x�y���l�����}��0���V�i��Q�ߧ �F4z��`aڣ�"p���2;�
	(�7��2���~;�لs�̥)4�X�,�M����H�}��Yt32��Hdg���0��O� ��\�u� ЩX� (s]�|~�O�����5�����t�b
CC����HJ�Z�ݩh���[Hf:h;U�`�A����vf�D:?a�=qZ\��T��ho�Ú����������L]���s�rN��U��'x��K�ϓ���U�F2῀͎�� 1;�E�c��{���ӗ��B�t�RaT���=���z�ϥG�睸��/��T��U�1sp�!��\�/)p���a}3�b"�za��Pķ��6�#J���Z
n��h'\���J{�q@�厛͸�l���q�٬�����!Ŷ���<��(�As�R��|��X_���]�ޱ��&L�Ў]3��\:EE��ޛl�c%�#"0��A�i�ɧ��
������GMJLN���\���: �M6Ӷ$(�=���ތG~��~�ȁ�#���K<���	�j���&3=��N��,E��V�����|��'�q�B��|�o�r�p�n��T1'=�3�y�}ݩg��#|�(Y?L_����V�T|i�b�Q�ۅ����۱j���� ]�����>�$<ʗ�3��c�'��Y �Q�l�3���ᕅ	�s�0���!�"���s]w�˟�Y�KzT[+ɜ�:C��������Ͳ�K5��.�*����M����d�����l�H!�ڮ?En�R�s8�E[
��ܜ�|4�P���8��I/ꅏ�m+?�����J�6��9wSUom�*E����&!
zE�DR��D$J5��e����q�hWø�௮�A�k�Ok������x�3�WJJ"�5�} �>a:�gAh֩x��}H6����Q.�����g.�7;<4sRQ�8YY��C���}��Dq#̤8`໳�����������`��^tE�����eډ�����=tV��~�&!�F'���+��RL���g��CԵ�����}�_��9�1���r8ĉ5e�9C�'㇩�#�~�jŋ����(l\�f�p�S=/XY��>Z�Dd&48^�I��~QN��R��1s��]A|8ɎZ�MN�#�L��<aex$4N�)�p�'�M�w��4h�O�dy)���<)ʿ��X��3�� ��׬��x�`�|�ww�+,+h"|"'8���mV*@�'��/�.�K�wb,i90.U���5�zP�n]�.�A2R���Fq�{��#�.e f(0R�${,�C	����w�Zڂ��=��S)!�II4(��{o�51���CYϡ&�A�����L)P'�D!��D&>U�P���Ҏ0��jCl���Ȉ~�����k��	�;n�4��A#���!9�&kJ�`�z��Olv�௒ln�\�1�Q>?3#� d�����ٍ2`8�O��\h����_@�ho
Z0�=�bǯ�1p���7�۾��ma0mm��w������Vd�[Z�\C�0�����[$B��7���N[;�YX������C��\.��{�:�HC��v��P
ˠ�7�$�S���n_@�~��t���k�	~��8����<��/�^J��kN���Q����	�:��ϲ��up�1�+�R�d���C`�u�n`^Δ�6�)�xI՜�SZ[W�Y5�*��LP��.��}��퍹�A�Q�Q:�c*'`! 	JNR,H�{�c��~��D���� �?�,k��;N�.����DL�1�J��Yk2*$F)ݿ�ŭ���?��l�*��@�2�P��t��Ov.�����7�O&���ܠW��0��YN�)�w��W�e[��6.O{�}k�J�	��(ᘉ��W�g��f�)G����U�/7�R�N��ot�}f�1���'�Q�(�����(�������L̅�oj)���d�����X�q�"�
(er%��[�TLշ�0��
�l�M'o�@�`'�f
̰U�6n�*8�g.�:������$�xy�x���ι�t�P�iz��H��q��'��Fg������#�M�4�/D���E���/
RE퉻���UNs�Ȕ7�I�Bڼ�e�D-"�����mXG�p�mͶ�U�]�fo�� Ǘ���X� ���%_庆9�W�v��0U�t6۲���?�r<�A]4J3gQ��ūጒ��J� �qɳ�K�������hx1��M�L�G�ۈ�PXn�Y˸Txv		br�.
Mݹ��w�/�bd_�i����2�,�Sw��Fj�'��aJH�<۲�3�x�<�h4��/��(��Z�B��a���Sr1%Ye�a�3C�kT������Ɍ2�ΚlX?��ލD��%�L��� �u�
��ϥ����t�����j}�ׄ��N�"�]��Vq}��h�zu'�y�mC;`1x�fJ#�����Q�I�t�cj��؛H�9����o�r{�`�d���H?��[�#���Ue� j�6�g2ĩ�-��eq�Vu�cjT�ƌy��IJw�^x���o=�ɧÔ�J�r���0��D�U�)�C��ͱ9V.��:�W�u �2ָ-�^_[�`�<W�|��q`�=� �>�y����
'%Ѿ�n�튁i�/��	 ��#�־��-`ِ�@v��#�t��$h0��y��D�J�I�2�2��_��X!�ֆd��*+����(�8W������ %�R&u�5��/�W��2����J���
X�~�l}p(/7�W��"]����p��6-�����X�}Q�^�5 2�ÆuM��i�\�V!y8��Jv�#� n��ғVo0��Ex�1��6y�u�r_����Yl�!el#���Qj�	QZYb�����q��3.�²��~ �ɍ`c�%P���<�%�v'*��'���0�BBC���*���@ϟP��:������ɣ)%�à8�a�+M5N��.%�&�����7�Fu���1|�=&�?Ud ։�8=X	��'��}|5���@aKihyeLfD��X�2����*��]��u��λ��}S�NJ́g�6��U�uv�8{� �S���z��j�'�Q���2h��2�<u�!ܩ�ʹK�����B;��>� >��5�ҴB	�l�oǳth}�_C|�x�������rE<,�G��·���\Q�{"b�o�}�\�OL����_������JV�6���<b����G����<h�9���5����&��� VZTM�h�ͦ��2+2;��&��ѪC ʍ��;�ჸ��J�5~�<o_�d������*��k־� d�[I�W�l�V9�m���U*6G�^�1`C+׭BuV�3�4L~�I�u�0�D��E#��\ Y�AOe��]�R[̑��=�=:�U_�U���l�z�X�i�ȍ/�v^Am���f�b�i�8j�,6�'���(�G�����5$�4����.٤��V�}�^^�"Dc��G�E��F�A��ҧ�!1�U�j��I�:[�SD��+���H���N�ܿ��5�y��WaJwD9VԾ���n6A��B��T�h�+U��4��7���~S��e$���%,�l[�x��gl��a�C�ǻ9��\��R:`���l:u�� 7P4�fC3������ھ�IY�mq������o�?�g@�A,z�V!�eZ�A���\��%.��k�,<ೢ-�t��h����/,���X`�FІ���^+�Z!Hz7�K�������i�#@��Sj�k�A[���^��U�V5�����n:r��aK�JjϚ��guT5�-H��<�u"!����xr�'�}�=_g�N?�|�vX!�F߂��{������*��l�g�.����w�� ����MCj}$�Ff����W-h�k��E��$���@ �>mip e�Yf�oA��=?��f�j��-y�|�F"|��/$�ޏr
E^t1�M]|#`�\,޸�v��c�s�Y����i�6�qx�w�%��af2,�V�m�%i�>f��������῭����ص6���Q�Jgv�V�%�#��o�o�<�b�S�|S3r1O��ϴxԣ�E0'�3M��@��8J�%O���Šv�#��$�mu�+wqv��^8긌�����#�
�==����4���{�h{�n�c�n� �����$ȶ�a1�C�?�'��{��~�1�r9����j4��o�e�������+ԁEG�!/��/a�o_^���*ԌHo�P��=�?����^�m'�[J���U,��^m��zV#�V�F�ᱩ��"����6���Ps7����%���B���@ VB�Ӷ��+�!V�eVΰ9�8���0M���*]NCK��"��䴔)t�6=v���4u�x��6-���ǆ���󉠢��i��`���r���Ї8��+fg3�
2fU-�v��e������Oy(���Fe�DL�DK�Sc��;��?A�����nwd5�1PeI�z<
��������p��wA�{��
&�ռ�ⵌ�hB�]��\��z��ܘ����I�1�F���7��~�^���(�~ö�#BE���ߜվ�R���E���lGt�������F��k���+4��l%�X�z�f|�
��/�,���	 x��m3%�ϟ���O��M�ް��
c���H/�e�r������F���L��VM��|:�������;�7��=�����ǒ����q!����j{das�n�b�Ἅ�����x\WH!���(���t��^��rb�s赋�~����|6�Ǡ��O��
�ڼ�����^f�H\쫆��U�Ȍ��uj�֚��~��SG�E���k�m���{��03�"�\�<9�����P!bA5UD�:�0�B���l�r�2r�M�Ut�>��k\�����j�F��tV^���>��	0��!����V!4�G�-ƖuZ�Ŝa�&s<�wi��&>/��;�T	ߝh��W6���A[��#4Q z� }�~��Mp�bpKYuHh�Uu������|ȣ�����м��(���ƓƸ+|�I���7c4����S���(_���NYf��4��r#_v!����Sk��;]�]NY���3�-Iذ�Z�̓O�~������3@iu��\�*C�=���q�EY��Պ��_��YE��Fo o�b��֖:���y�KW^����/�E7�ˀ��J咘��Y�P��F���cɭ,���}a?�HGHX�n�lȑ��勨\V�,��j�l��.�dʴt��L�';�BV��������8MjWR���t�m���A�]D=0���㨉�2��#�Z���K�ӡRQfY0�jbR�	A�є�1��)������`s�G���ネ���֦;�ft��1���!̞C+b�=�ގ���[To�xH��б��F���S��`�
�2���0�$W���=�����@ee�m�t#�:t�+7i�k����a����x��{�u�8i,��3�(L�Bn,��+���P��J�-�+�C;Q@�+s�z�>Ժi��඗aн��w��n��oo;8	��(�����T���`�՘�%��������^a�C�Q��8w�~g��#ʜv�io�t�+��yo> D �����������`0�~�����¦����[��u���I>T�A�{T��8�h��K(P?v~�50��?Ig^�� �d�*z=�	��X3):Q_��8y���&�%U�ʕ@2M~��6���Ϩ�G�:�]|[x�b���УR+�5�<�JF�rמ�F���t�H���w4t%�nؚ�D��K�jV� �MaƱ��|�Z�B����T�g�qP�h�-M��<U�P�`;dv�`��SC���'�� �:wѥ���1UMc����"����=����H��|н���^iy�]�'�g�uc�e��I_E�@��εeC���u�z�M�6]��w^l��j���Ѯ��U�f�+r�k�9)�j[���:d�����|�R}>����>8v)�yr��r�I�_��Z�"�ūP�
$i���!0$+&��~����̖1�Fh���́'"�m �$���\3����7}%*�>��������y��$GՀ!��f�e���e ��.�8h��}P�N�J�����z��'��Z�vK�{g��yF�^�*�wh�G5e`wK�"Oʗ��]I18^��e�Z��7b=�;�|4d� 55�f6�v���eQ%�+��o���eR:��	a�s��|Uة�h�eI��8��bi�	@⦝rޜ��L̂ds���Uzӯ���Zc�噟P�5_7�gi�D��o��&��_%�=:0��E��L���Ch�9���բ�Xk��h�H����lW�%qK�Hnq��y���fjH�;ęg������ˋ:5���F�b���}[��;l��J"�JX����!q7A��c[lCq�V&M F{Db�GG_���6����Pp��c��J�6���*���n��f�S(ڀ���?�P��C�y-��φ��F�9�7 Q�[&�e����vV8a���H�<!��ġ��*pg([�צ%v�ʑf�b���K
�k�>��^�)�xP�b���10�W����y4���S�df�/|q�t	R�Ҷ�wۨ�V�&�7pPjP�t�|�TN����E��"p�}�Ԯ��ʊ�oد�4�7_h�GC�Գ�Ձtc?:��֘˓�F�#�oԡ�3W�"?��K@�˝.u}�2s��>��G�����(�duI<�:�
h;�����%T���@D݇M���
!��5z���Ƞfe��Q�]�3��%��	_��댘�4N��AE��2��Cׅ�!��d�Z�}͑F����9��{�m�}Dm>3hU?l���o���g�ȫ���	W�锾�XZ��H	By���x�r(�$�45P9x�I����L�S��Щ�SR��[����#m<���j�lT��!CjKU�|���1q}Զd{�mݭ#����CI�W��>�HlQ�����wq�1��@7����50�����{*TqkJ%���:()�b����N�?�P��T|��?N.�9�]��m�l��$�����wn�Ӕs3�f�c|f�/��7}D�-��%����۽�gE<���+�!�Z*�aT����9�_zvf�Ot9�iW �LH��}-�㯉�RM��S��'�CR����K}Ȟ��\<qd��%�u��M�XZW>ẅ���l4ڙ�ް{�ѐ��<R���=�T�
A3�+�B����k�� 3��ӓ��Ρ"�� ���Y�E�݆, �냻ȡj5ֳ�?���q�~7!�?]�r
L��$5�]���%T�GE��2����4oN-_�Y�s�Mn��2^Y�::O���Mu�(�q��](�am�<x �;�Y@�z ���^�\�H��U���G_�������K2#O�_Q\�v�3�����ʒ ��Ʋ���՞Č_�Z�A �u��H"$S�[/�G�c��V�a�^�WƢ��Z/�H��_˺�)�E2mAR1����h���[6����H�=_��NpU�\�"=�!jK���=i?y��zC���͇�}�2w��޷���Ni�)��Z8p;bS9<#h5�T&b�+��2w�8܄���h�������Kf���bi���^~;
�����Yb�����74d�5S��LƲ��o��"nv@�c��V��HH;ޱ`"G��3kڂ(g"�Oɔ՞�	�l��A~@Py�^J~E�0 �������zz�����T��%���d��|d~�\��@���m-a��)̄��濾�,��Cq� 0�8.T�^;�~0P�C����t��[��4��އiTl&��ǂ���/��%I�Cן�
��礌QЫ��kQ�=6
:���;w	D�.��&>��E��Į�N�����9��ï4�yTn����[�����w*��kr_d��c�8�J�:�6�ev������l7�a�N��"�`ƶ.�w[�I����,��!�^�W##�$��ď�O}���'0���7�����"��������9��E2EʪK�C�	)Zv}^�t�֥e������͵�1#�:��ôf�=�w�MY��}�r�_�X�ȔL��f{���BjmtB�[�0j7k5a��+\s��ݗ��+�C��$�EQ�	�\D>�K�;�a6e��b����8d^��U��C����]��{ј�ěx����_�Ҍ�1.W�3M�6��O���{��愔d=l{=�6��Y�rm�Xvx�;��ࠕb�&��lP99�b����}��f�aH8���0�
t�o��m!L~rKbAwo��\a4��ݝ�z���C�s��_�0�i�I?�ǭQ��kV��2�v�sF�.ؒ�f���&��{"�	��?� �l�\߅��9uX0!��;ݝJqѳB��:ǽ� �X�k�����5B?�B�ɔ�`A��f1���K_�Tq]6�Ӈ9� ��.�ϸ¬���5B�b��ǡ����+?��4�{�ԟ"*��=�Y���wC,��N��l0�����%������B��N�G�����}yp��������Tu���%5�b틓s=�8;z���?������Ub��"����"�j�m{%�zb��fƞG�	]f�k����)C[Xg�v)Z=N�*�l~�k�	/*?�r��?��0r��U�ց��s]�������}��-DY�5��8
��*�m6���:���c�,��{�p�X�6����G�	4uRb�C�T����R�c��㕔����=g��%g�ស5�o��@F��ȳ8�\S�Ԝ���W�N�s�� �A"��^�s�.�Krv�4��w����e܃a��d�����f��4���)�|%o3JϤb�s1	�S� ϥ���|Q�"��ʂ;쵣uq;�2*e�炮on#U7����;�s�Nj�m5-	�)n�!�j��:D�jtW���'��Ω�2�"q$�^}'/�>ٳ�%b�n#������+�ZO�5����<��M��W�6S�&�w%��.�>�[4KO� �����dO˙�
Z��K�Ԁq#y�,�Ψ�_���6`����݄�,\��j�M���I�x��T
1�ˢ����e&�s�������"e!mM�v���j
@}C��yG	]��O1h��e�%�d�-z�BEa�@�^�]*xڗ�Ҷx���s��W����y��O���7��(��Q��u�#�>��ngU�*gYΪ~qDd���Ԅ�i(jE �/��OhT�;��OM�B�u6�"�͇;(�W��B:|��d4q�������((!���`$2�F!B�>���+.fܾ��gW�Մ�3���P�+�lzf�aA̺�-M���U��3����N���V���=�� �@����%5R"��s鯩M�j�vU���<$�\�������LP��
�N��%���6����f%�F؊J�@)mz'�DN��w}�#)@��:]q��G���;�i&��d������ c$�*!��8�T��kV5�R�\�ރW�h��R�Mo�J>���I�Ц�fȿF)m��&���l�e�z�%�>��o~���^N)����!�8��rٙw����d��ZL����:�k��b����T�.���0�S�- ��:巯�$��u�瓋��͓c<���,+��b�Z�\��9�5��
 z\R��81�!�q)��+�O�r�����Jذ��Mi��pՉ��"��Q�d��8��*�{M�P �{l�u2lz(�$�����
�U-����-�com�Z��� 	��y�⣠Y�a�1�)��h*�tG���:īĳ�5bI��S���>8A�ӗ�I��
z���ѱ/E]��5�hSr���?�7[�Iu�n�P2�r�n, �!�BB�D?�R����"��OiahgН6�鎹ͤ����~>G�ڳ%���$v_ }n�y�wx�Ha"�9���AC�󳹔��qVnk���u��v��΄$�޳X4�@hNLV.����������	S�L:?�L�ׅu���x���@���$yk5o����679-��_�l��pB�ܷ�喗!bǂn/�4��=/�x��(��x�bK���w-J-�m��
 ��g��m�4tG�J���{��ҝ���7e�F�C0XÚ�~W��:,�����@��u��Ml��ޏ�.x����R`��B5E�.�S�	�:��0��H�E�n�u�IЎ���sRK?i7�xCS3���-��X�bPY�j �h����v	_�p�nAvbt�mQݡ��K�T>�R�U���ׁ���T�)rNQo;AhA�c'���ψ9��f s����<7��K$h��k\����;Ü�z�:��ZS�2�I��A�loQ���]�j aĕV�z|��@%�-4l��2(���@mN�T���dN�� �[�˸?��'�_�5��ݱ�cH�\�p�EY�Pr[��'�G1�#�sk�W���U��/W��S��V5#���"1ds��s�y ��w���$�e\�T��MzZ��7�GvR�Ռ�Ad��`�ag��)��Ȝ}'�U�YD~V��z[g�,����汄�I�	_^��-܄���T\��h��#��~\�=����T9g�?�IZ�5|���w6�Ƨ��j�֦������޺/*�>_���%D� ��.��qp?�k�~7X{��Q�	���`f��_���/������Y���@f^;q���|����B�1��6��X��T�WO��1
����U��2c:��u��ĥD��B�-��3����ī�PFP����KG���L�^��7����������U�q� ki����i�ӕ���n-���A�(�v��_ҥ
������C�mCt��,��|�OU̾g +��"�_@@������f�rEֺ�p���􋸞�:AhB4ie��䅵�Y�r�3��t,�ןr%?~��O��R�bf��2bl���TI�)����m����]��Z"�,�B�4�\�����o���>�4�����-H��:7��6�M�X~��I�$G9�d���*� 4��;�0Ί��<�=~2�\_�{6;վ�}���c`��p����I�}�>-zͷ�8�.��w��<���f�H�Ҕ[��d%���K��]U��UZ=*���e�?${J��JY����V�z��1>E��}�::l} �����]>7�o��(	sN�����$�m��*L�'�x��v�wⰖ�P.��M���;{�A}F^ٳ�Y���� 0	�K|���1�q��!�&K�@�S�]�iA:�����bq��8-��7��Q{Z!A�X�dH-'�������$1եc�U6��]�T�w�IT��7^
Psx���X����x�b�F�Oi�bT�H��妑�!�S�y�e�3¤q��P�K��s;�B�_�C�R����E����,�5>t�2"�9s��l���4�.�ߢ\{ML�%ɫ�9PM!���T9��*�7x�ۿl�Ҟ�����8p0&9�)@����~��<�1�U!)�0���d0�Y ��AvR��7V��;lYq`B����[��Y]\�
ŷ�/d~h�zLe陈��M���]T��[�0�~��?z=�����6�#��zxC����Lh�Cl;}���О\$�]�?��+|�Sk��k>�H|A�����H B}k�m��
���-����t��w�EYץ�S6B�}��fð�K Xaw_��9T$�׆��W6�Ė�P~���8qNA������K�1nA��_N,�Z"T��r���*Y���4���;��|JG���˖1OSxA��qy���?��sǐ�^��Ò	�-;��R��2&s@��c	݌�-4=K�+�l1[�Hc�_�viEiaB�7��A�~I�r6S�V�'In��2'�l�O�j�eH�lh��H ߱�8��R�̕`�~'���@�4q���eAF���LK���q��t���@�I�@��>0A�������@j���p'����2,�g�GW��{܄'u���O���׿��mfF��~��'`S������c_��@�m�8���a̡���C�L�%0U�|���7�w�]A[t��S�i�E�4~4{������h[�E��0�BF��]�����O��q��+�D���]�v��bhe������J��N~���T�pn�n�W���ğT�n �<<�;V;�
$�]�+ �%��� ��.��݊'{�Ҳ�������M��].��R~�9���1�pݩJ�F�g�KU���,/y7����9p����S!�!T��p��|�?�'~�hy��2�TI�[5��F}G�(x�=u�ba)hUZ���`cdr�J'���DEyc�U������x��lP�G�
q��i��TL(Oc2�~p�aOJ�حSn	F�^5h�N�<�.���.��@�b��/v?�ـ��*[I�N)�� �w���q?#��ۼ
�̄w/����d� =�Y>��6(4���3Խ�P�bxA�!�K$��+�h"�A����xe[��\�Ho��*�-��V��	K	�7��z/m��^��|��t��_~���`�w]ޑ=Q�fm��rK��)�AbW�
�M�a�g����_H��ߓ��E�a �X�ݢ~��>��q��|�j��M����o��ﰛ�����;@¼�.x��C�n��X��@D�7�˒�-M^�t:O���V�����#,u���⽧��%ǫ��1�kV_˒<H���[=�$hR���\�X�U ������KQ��~C��]�R���D��MQ��<�v���q{J���j�!'%��j[k�§`���xEO�I��J^1�2�;�G��>��Y�b����q�jj''A�9׻��j�h��J��,0�7�c�!���P�D�e�>6o㚤�к�A�)L.F��|�@����o� ��g�,X�loH9[�$�����,�ƣ��D�i�ݕ��O��C92}tB��a��)�AN��6_s6��ϫ��X�٥�	�њ������8��!T�0�*:��w��n��ȫi�7WO@�c��"s��i���m�dR����L�����Mk�K:X�T^Sb�6!`��r��5Ib��aǘ���租3����Àr��)�h]�X^����~ޫ�t1e��x0_Ȉ�պ����Js߻A&���9�pZ!�8�~`8����^��6��H����"�]���ݜЇ����_q� #M����j̘70�9�@�02N/���?L�,���������񰈛���jTח`x��!�_���R*<��d#�����c�&�g�tϏE2YaD�j���ST}���#����ohqO�hH%S�\zԪh� ��Y�>�jჄ}��g�����!h�R�����O]��y�=R���Ns��^DF%7��d交������5��"��^�!-?"%jkԾM�<< �E�J�"��:����M��\��(H���lG����Bg#�
�+g�������|A�K^�C��k�L���(�_�I�JmF'���w'$����c[�ϙ�hq!������\z�$Վ�%~� ��`�Z9�'��w[7����cO����6t�s�J����3���O�'$�K���	��>4�h�,��~�	'WP���O���޸�/"6��P8t_8"֩�l�i�,N�2Fd��49�ͻ��cWT"ӟ�_g�v�kE���h�o'�K�X�붸U'�\6��X��q������*&sp^�C�Uq�����B ]��8���В(�"�܊���J���9�?q�:-_�9x��6���_1�h~S��jc��]���ԪC��>�W�M9��ȄYb�Xp����m�q609&�wHQ�O�S�֓p:x�s�W�l�J���wlP�%Ƭ��˟�A�YJ���"��?u���q2h&�&��;��Y�;o\1}���WĽ����Й9R$Aiv�Kl�I)�'��L�)���XXO�u�s%'wzÆ+�҈X
�}�n�gP\A/��L��&/A/:C'f_'K6�"��N6J9MP&n��&0�����J	��a���^��\ZqK�ϕ�_�~�(��鍶��e%����l�S��~KA���|ڲ|���;-�)$����uA*�x'�U��7���$���'���`�������m�tM��V���[����b�rQ���b+�<�k/qt"7���UM)~32Gf,�n��+B�� ͐�*���ug����~�3��#�
�������O	�N}L�(SG7��v`�ˏ3�7Mes�%wF��o���6��&�ʦ�奀7�"΃���{�87`�?�~TM�.�C��П�O�QޯH,��@�˶�.����ǦL�,D;x'��.�VGN1���F�4�N;�.���X�1����C�">n����9���M��=Iy?������g���DA�V&�L!�4�W����N�,�oe����H�҅z��x��Av}mG�v��R��`D:���e�NȜ�$���ò�&i��ٳ$M�z�$���t�@�;Z�g��uU�m9:@�S�hB��1��Vf8�_@�ee	;�Fs4�;��u���6��wX��ݯ��z��<���RLa�߭t���D���U1��k�B�aF5F��9��?&Nt L���Ēӳ��%ǉ��!��q�K����{�iq���o��wq����s��&��.��L��y%=�f��C:/�=/�z�ε8����x\޿�رj-����.*�\��$�����VP�!�+��T�C9E�%��& ��D�`	~W����B�u(�l�2C�9�tS��������Ƚ�H��Ǳe�����6� ]���TԮY���>��2�s߱í��!��`�,�K3�D�$���X��Nh���S%=�:�ii���еϷ��"%\^���(
m��Ŵ'	s)�'�)�8����~��
�h�M\�/P1߀ύ�b����]i �x$��`�ڣa�m_5�2HD�hu�g2��x�Цd�wt�r�XY��+"��)V��O��e �������L�Rre&���]T+\a/�WڰH�E YC�v~9K���/��x�3�;�N�G�M�"�ٰ�����|�J=s�Mv{��uI�
���2�q�I.Я��w��oFU�lVC���𽶬ܻ�/;I��n�DίԔ8?c��_1l���F�ַ�����-���!b��1-�L���sdH�i���d����@�x�0gjte�k�� �B���}���w�J��^1'H��=$�j͋�p�7�5��UL�l�	s2�:�� �����ق���ri��faRG�f}yÝ��5�Ǯ;M����Z�
?����*�x�Oc���_�L��gc@>��48'ψ�o؀4ߣ6l�@6h�)��Wڠ�j�5=���SK>�΃�<%S���K�o���GL�N����w�EY�9����A�wJ.�pe�u�ۿ�KS9�5��v���S��B���Q�E^PW�R��+pvD�kfH���q&G ;���hR��M��7s�wP�
���Y�Ez;�͒5`�w>=|�h6,v"����ْ��Y9}=zU�<��T�2ј�\�
���Js~7�H�_3��E��Al&���,T��}�YY�A��
Q�����crV��&�q�-��(���
�dU@G�&�|�b�!��F%�KX�.`|l�-�5��L�Z�n
����[��zح3O��KxnM���f�<)�����ۀC�4���z �16@��#�?��D:��Gb�u�w���{�IFg���>n5�Z�(]�t
	ASJ��N�!c�X����l"�R�D�T��j�(�V'��j�$w��������j��k�U	��Bn\��*���<�	n�����>��k�Rҭ֥/'��� �K|��.�A��׋���C��#&Jka-u�w���(} k�/{wN��J��1J�n�)a�C�!c0'8�p�/َ�
�~X����G�b�ގM�Q��v�a���Y�;���{߀ �i�Τ �����F��wn �O8�� ��]��Vi�[�Y����= �u�֘(&H� h�lr��]tb�?��Z6f>�v���sxӝ�O�R�����y�x˯����/� Tk <�a�τ�r�rn	��Hb�)�u�o�rf����cz��N�i�*c��_�@<�䀄���z�O��؏�&;>�>����\��>�O�l��*V���2ʋ�s��3L���;�a���-S�u����x����2I�d�=�3w��9�ȰB ��Q�TZ]�bQ}#�5��A�u%�ؔ���pT�m&�clY�S����z���|�,Oe2�Z�A�����,��U��\���nq�+���ߜ���A�<��`�_M�,�a�$�'���_KT���{*�>�����#�Zғ��[�����<��A�d����SaK�ބ�*Yk�ރ�@��!w��-,�>�_o52��|M�Ǟ��6ͦ���HM�'J�5�He��80ҞMaB�%B�mdzc��;���p:f��?'�͉��RS#�]�Si%����N0,bUK3��+���v�ԧ̮Ē㪦r��6L �
�.���N���� .-G�h$�	m7�"���
��~��0��.۸�$�)r�-q�)��F��SU�&Q	&}'���&� ]�Ò����[���u�5X�s�����wV���F(���Drd�?C���XMy�FI��E6fsP��3���jY��N��:��Y���&�$�c?����59��@jh��t�Z�F��q�@b��3���_�DS}���g<�bR�˯\9��g6�!�"����Gn�%��{�F`/IV�����w��q���Ys�w0�.���5��OV&�b���O �ӚZ~�Ae>w�����rC8�� ��$p��y�����L3;m�����'g��Ƿ�<S��}�� �U�'�[������DQЈ�=5����:|M҃��=D_>��=�6~���%(���0�eR���1���L�,�j�c*��}�Z�?��t�U ���6	r��vK�b�A���D�x=� ����z����P�%޽��<�"�������6�Wj����D��������AQ%���5J��E־���s;ֱH�����{���an�;�)�Jq�W��0ӃWa� ���������5�%��+Y�8�ژ�a��Tl./��?�+;_􇞸�j]�2]�VD�W�o�$
�0�I�(m��*�M�ߪ{O�=q�,� 9�y�X�,�|�!J?��s��g�@p�WW��Lܴ�Z��'�๺boh�a�l��"(��=��F��.�D�'�u�3�yXס�C���
���W��e�X�Lµ*9�Vrdd}^.�Kf��ߓ:��
��X�W�?��(���
G]d ��p?�1�~�Nk����U�􏊁��f;���9$ˑ!EO!.])�"p�9��:*�F�*�EK�N@�4(A`���W�F����d��?r/�%�9���g�WhSa�������\�V�$�K.�bp)E�]�̂��S5e�h�)a�������/6i�l��΢����Xs�3��\���Q��^y]]Ķ.D���[�-�JGUܑ� ���9X׷�E��:�$d'�!�D�tܤwC�F�-#2�Rq��m�7a�6~��Q�U!BJwU��#����!�'U]3�^'���$�ZM�S���"=��SJ���%㧧�
��J�C�y�<D�zG�,۹TJr8/�f�>�h
-��M��z���Ni�@�o�w��&�*t'^½�75�U�=gL�y��	�')"�l@�>^�
��dd�Qkt��_W>�#�y���Dݤ�-QF�Q9Z�*��
I����C[}���'_��d�����.�.3'u�&��Ii���"]\�}��D����y?3�t%���̜j�G����y�H�@���!��?#�����r�Ȗ�?����!-�a#�^R:Z�t#*g�"��[�,'<�=G]5�W�3:K�8�e�k�b"�ԛn*o�E=0��gf�3�L��AHf�%���r*#88�m�Vbm-G�@�|]{���p�hȷ�H0P�ޖ�|Ժu����>M�{Lq�)̒0b�i�� Ta�^���g��ه��j�U�Uv����Բ�'&~O�W��IZ;d�D��K��ˠxpR���sK���-�S�:Ep���+g�C���-�H����x�5���jQ���dz�;2Lh5�-�ƋU��yAI����#�E���4��\^�"0AR�������W��L�| ?$zG�%lƖ�
Rv"��}������}q�85|ܳo�a����Iea���WD!l;z����pW�Rq�OFY�
���:��˅�b�q�*��Ɋ��cub���*�臅fS;F�mɩqdi+�_��U�Q�'���%��T)#�n��Xr���c����^�qZo����4!�w���:>����@�SXZI�����F��r~!C-I�� �<��S��b�K'MY�h���h��ͣ���r���C�<5���F�k�[
 �nx�0��J��p���B��
:hT{SNiU��X���Zo���!,Z������&hn��������2ҝ8\�j�pGҔa݇K?� � ��|��;h����TdŬc��zi&e�2�=�wC�K?|������]���c&0G��XL�T^9K��a��i�X�C�|8t�M�PE��[�D��U%I�����@>�w|�7%��{2"Z�p%��/A�L&c=Q;�S��@��RI�����m���,`�>�����@P�+=ǅ�� u*��?�D?��U�Ǽʄ��_.|;K{�$�L�觌�u'�P��f�kܻ~��U��F̄��%\"���o���D ��M&=YUW�^��q�l��_�b���>�;��aF�Q�0�C���Ub�4��F0r�C��0�ۍ���<�׆6�9��Q��w��hv�j�oC��y����H�����(�O`�O�8�2�:�yf������MWh�?�&@x`7���](2D'�e��P��|��~^\o���<���1+��b�\�uB�B}����My���� t������M|���}�1��,�K�?�����<^X��d������~�K���%�O\��!�>�����n/����.I+֨�Nhҋ-tq��E�B�xcL��y��2�������xoF�(����U�3��eq�%:X�	C����>�zbSE��Y[�p�i1w����{�@�~� �u|C�q���*ٶ�7h46�yNtk����=okoZ{�^DV
�y#]�l��&����a��ړh	Y$@4�f$f-�!��o�\��CC��Z�ƨ�t���zJ�<\\��߿�̥�c�T`�nL�ƪj�BE��4)�""��$E�`��i�^�i���rx+�᩟Yr��x���T���p"�;�F/���(>�$ҮG|슽:�hU�Ov���ؐŚ܍f9'xi�`��)V�J�IJ ����T��=����W��Z��q���ԡ}���j���j;.�מ%�A�B{�qt4���2�N��b������1�������ǘ�M�#�&G�Q]ck3�ٕ�=���pn�7��G�R��B0��x��P�+B=���#*�
����H�8[%�4z
�b@���i���.��$��0��S�1��j}c@��4~HY�s@�:����:�ͧ�Ӓ\AN�$e��m���/�����=n,��kȓ{�D���B�؊�f�� �09�[����8�l���k����U�N�s������@���0C��~��*�Z��Mo�OW���x���ϳ෯�^m���y����e�	��P�T��ْ��Z
m�g7���B�4�+r�m�Bn�i�ӗ�8S�E�$�S�R�F���PZ7�D=���P��<�jZ+�(d��1�!��G�0=b���q��Z4��<���`��XЁ��6�=�Uκ4M7���\�_X�5�utU=��/zXɀD9w�@7��A
��'��ªF��QN/w|�S&z�)���9�l(��vɜ�3��s;կ�(4 �"BޑK���v���6}�&�k��0y���d��J�?�ʼrs͊��qm66�?NW�	I�1j���	����hm���Vy�6X��y�
'Y���ۓ��N��Y=l�G|�B�B
2��:ƭI�\�'���^�i�n�6���=.A�,��P.㩵��[l�؎�5˨A˘�x���m��9�k4`�]-B�-lm��C����[�a��Ǆ�%���W��M26���+*�R�j�p�;7n$Cq�L�8 oo�M�V&�xX��dڲ<��|@�]�^Z7���e]�hi&�j%}i�AZ� :��t�j�Q��L�3LZ=�2#�0&���S��qq@)�
Ə3�dVyP�Ͼ�E�rQ����<��X���S�%EXg�ꂦmmPm�����&�_�,m��(
�5kj��v�,���3,Z�,�TX���U"�֕�9+��H\vu�t֚��QJf�U�3m�s%},M!�ʋ9c���͒k�����U!�8�:c0\�U��`u��X-�"���,%"��S��	 ��5���'CQS���`��z	&;8��$ݡӨ+^��G�62GQv��u'#�3����$�a̢����6�@���(x�Y�08mǨM$�������ή�	�кV��;W@�z�tJa�0`G}�]x�N�9M�����q��\p*�8���_�WFc;T'��2��Rg�8L��ȸ�(z����f�XK�����v3��}��9���ƌ��=D9u��z��`=h2��P�KO����6�����!*A�}H)�0-�	v�e�F�a�����:��9H9��3����u]<g#7�,&�@#ȁ�S'M9;�(���C`3T��!�V�r���;��&�[e0O��+&�7��_�Ϩ�I�7_$s��|���� ˇ�ɐ�	CW�rN�}DHzmI���5�$#=����3�3���Ey��)��~�?�Ш�v�'>p�6v��L��SN_�l#�����n��xa*��3��syƹ�S��|�?H��6g=;5浉[��:.t��sL�yJ3'�kB�}'/[�;0�\@��gg?]9nn�xr?�Y ��{���Zm�#�1�	]�o�\�p>IGB�Ŵ��$�Gb:1���24�[K�����mq]��lq,������5�A��0�c�RCG���/��#��(�֯����%������Y]W�u4u���v"�$�Bq�k�dB^�bu_�y6S+�A:0?KUd7�sE0�9�ppR���2�H�@�����G4Y��#��8[�R[�&��ÀWbe��@����L�,_#� ��og{K���b�K��§�>hwA��bJ�5���o�p�2?�`&�d�ٸ�g>�Śb��$��=p�cC��	��RD�	��dk �IXёR=r�͘_�c w�ͦ%�~��{\eI9������͆�r��vJ����W�#�q0����vs���(�o-��ZElm����}�������zY<+ud��X�Lf��7� �-��L X|���2�I��x%�,}�����*�r%���9	[�G����BI�����f�~_ޕjU�m'v�.[)�E�pB�i�I���
نY�>X���J�>5^�'+��m�!�X���+��o`F6��TS�h�ߑ���b��[78FN�Ŧ'A��9A�]�'���'�`6B8f�<ӹ�)�D��M�b�P�� ��/��ϭ�٦�d!�G�S2�%��d���ӫ��ď{S�b6󅯶Xy���,�ͷ���U*u�fm��F�f��m�]�A$8�Z|g��P,)�~�+�u��Ы��X�*d����ݘ��3~q���1gy�͋�;n�Pڏ���f��� iQ��cdY��5e�ϛ�?Z�;ȍVzo����fTsz� �m�;�n�M?o�G������_�{�'�~ x�XXJ��,9eSS�.�lr)���J�@j�n�2�� ����H����s�vk����䢳�Ǜ��/d�\+��}�~��מ�VԪ |���������F�o�c>�;��hb��Z̟�;�S�Ҵ�0�~�GpK��ݘpm0ɰ���[��Hi8�%@�V�7ϊq�����h+�XT�t�L�6�#ő���[I7Ƚ�["hi�����g	S�P�ވ`�˝�|e2z�U�Wvอs���c�y�hB�ڥQKBȼI "����n�6�a�y�$��T�~����'���a��H�H:A��х����<&ϭJ�%<��
W�`�<��,^5��zH�J�螨�q�l����4�߀�>m��+��A�y������X��F��y�]Q�D��S����o#���9"e-OoЎ��t���,����<v�����#P��a�#��%��k��(ٟ�ٹ��	Lo�?�j�3%���q�,꿴�C:zV�0�AqO��w��v��@�C8�-�}����a�)H�
ݽ��MN�H��l;��p]R·���(�Cޤ�|6��p'�.:����"u���U�YM׈K0#3��Iغ�'�Wz�D�@R��	Ά{Q�1�+g�R��r�X�y\��;���d���#���"�ӐI���b�Σ�����Q�uL���ӆ{;'����x�Z�a(�G�K2:N
�!��ܒ!�{�SB���Hn'l���g^%@Lǧ?����WEv!<��1�z�E���ŨG��,�`D��0u�a}ټf\���.�N��W��ڃ$Y^\<�@���<��h]��N	�:۱���Ĥ+"i���݉Qw2�l��́������J���b�EYN (��p�H׾̥���>)%W޺�����-�-lkk� !�v���@厂ę�=�eQ���@�t�Y�� �[�y��]8fd]C�����/�#��������W��U�������G����$�ï��?\4�b%��~guVUB��t`��t�����_/k�k�>��}Ts�Z��z�p��O|�"�~"�)�]|�dKegS�HZ���g"7X<�T9�hQ<������ K�\<�#�kN�x\~�&?i�tP�R��4>����Ƽ��9��
RXb���5���,]�"h��(�DFi������}Y�b�!�TI������E�%�k���1z;'�/���"$s��7=R"����ac>WI{����������(]�E�y�N?��#�O�0"��,o4I��砉8�N�C�I�l��p��+w�t%�:�Z�!�ƫC�R���%*�.a�I�(��ѿ����W���M���zV��j)�v~���c០%2�2vIʡ�T���`�����$2���}_W����h+��7��|���*of�Qa���:�E���ꮫ�������u�wִ�(8xz�_���dx{M��v@^���w��ʶ^[������s�?v�oz)<0�A�-xE+4����.A��$�r#j�i�9��e���Civ5���P!&xK��ŝ�fk+u	K�os�FX
�<L"�H���#!�_�߅9S_��5��2{��CjMM�#�
��5�m�aJ5ߤ3�u�-E�����w�f@#X
�J�9s�G�`�",#tR�6�*�ܳ�f�,���~O*è�0>ʡ����=�`��.�DCyd��2�S�:�H��4��@��r2Y�����O�2���~Ǟ�T�[rR����of9h$��ᐪq2��CA��Qu`+*x��9/��W�ִ\�Z}��㡊P��I"$g������6�&�hq����DF�Z��nP��tm��O ����������"�r_���~�5�ŉ�F�%#\;�<2ゲ�H[�#,h�E�1@x����&MH��'�V��̾�?��Z������y���·	��Ň�;7C��������o�	-�Qc��Q_H�i��pu#j7"ao��~�?� �d6�+��w&�$�k5�]�!�%��b#!rL�P������-��0z�F�$uHe)�Do������inD�&s`�o���mP�M�e��S��; ���2�E.T6ٟ��K���,r��*Q��lxW�/��z��Z!ST���6�}I�~ۍ|,Us�X�/c��*L�4����j�?��ܜ�:�q�[v��LE�L�';��⟘�t�����{���w��ǵ���G>��>��;��?���s������gg�J�����]����Ý�����n�VP��0^K��c��{�w��"
y"���<�':��e�~$��@��^�x���}n(�
��RJ�fj�������2�L�c��b*0�����mP�`�N�Fd��|�ڊ�:�or'�h���8\;����ǚ�WX�T�?�)��sg�/W,�`l�=�#���w)�mJ�˷�r�Pr���iD$��ʂ�o8_A ߂TV���ŉ�"���R���<Z��}@8Ʊ����o$ iv�-*u%v�7tX��+��[�͂&!_�wKބ�5\��$�o��"d�++��,ڞk*�q#7w�A��b�	��8�?��PzpD��9rȻ���.P4�_ oD���� ���:(۴���IG��_�s��|����A�.�A�(M�"L@XC)6x�ܭ�x��t%�v�{\\�ek_ߡ�f-,�ċ�"&x��+Z�ߐݣ��b��7s��FnɸC�A
&�.�OW�^�K��#?� r��v�
ٸ��c�����>�E~�}����q=��J$B�����lX�Ccò�R��I��v��Ӛ0.�W_��Z�"�'��y�kW1F�;j���
���iy�D�3�i����}K�>0�]�2��ǖ�}��(̠�m��i;�fCiij@�L{�p��rSW}k
��(DQoi6'�kNH�����G��W���"��i���Q���<�K�(-=]�Q	�u��Fph0��/oES�����&b�	��p�w��"��rv��e�-���d=�����&��b8ş% ab���Nw�'e���\Z��m5&8�������Q�+��mJdyIz��vN��z��֊�d�`�����{����дK�e��X�Ȟr����{�L��
�U�OH;���HJR�k��n���!����ʾ��c���!,<��LzY=/Y�A�
�g�2T�+5h� C2�\�V��C ��9����w��"�w g��f~<�A
7��XK��U*i��E��1�B飘�hpQ���?�p�I��m�����T�h�kP�ƽ�{FwU�:�]�f6&����'v�8����^I��&��w�v�.����n;�i��^���L�������8T
V\%n[wBm�	x�HI�۹������ў=��*���Z�`�z�J�^��=�˩EoU�]����n!S���.�fZ(��0'Ͽ�������z���dIU�{����M�jn�cJy�!�Wq��^��X�wQ������)��!�ܑ��}>��0��� �v+2>�T����l,!O�=�tt*����`��~��Q����W��lY �W�(��5�FT�Ơx:R�*s�W��_��w**a����)��>�I�� n>�5�1�8��Q�}�����.	I�ʢG �?����Pt!&'�Z\�hm`�נ�&]��޻�8˟,Opd�;�1ɓ�p�n��|� a �w����f���~̭�mMNS[�"5�@�Ҫ�T�����l+/"/>D3�1�P~��m���Ų& �a�\����O��ަQf�6Ȥp��9�8����ӈ���7��}u̬��'�*_Jw���3�9��})�;����M�d�*H2
���0r�Mb��]�L�
\讂SP!eg��QQ9vG�;�����tRY�8:��aO~6�\D7�� ]BX9p�Ȯz#�+����gg=�쇟���P�0��!�������Ъ���-�!��r���稺ؖш�=j�W�n��ܢ�N�
���8�+di)���?�O�_m9.����/�u���j��6�Î9��2P��-7_����bn�,�� ����&I3����⺎劓S3m`ܖ������xi�ss����G���+m:��˵�y�����/ڗ���8��B �4Xy��m�j�PvB'Гº�c�֩І�iG��Np�U�̀3zLqa�ά�'���|L_D�Cw3ɏ¦]�7�>��G>F��,8m�e�%��h`��%��Hc����
!jr��I唚6��3���C�}.n�Q�5��� _%ȼ@�y��޾�!O!CpB��-{�����zYޤ�KP�#��<���sf)�MJ���{�*!n�7������#�.���7�?�g��|*���k����%�^� �^�${�#��^IY�^B$bX��R~�&�bv}��+y���Y��:�5�&�4N��L��h��F�~A�2t���Ey>`�S�f�����2���߆&� ��Y���}�ؕ��%��a6s�UJBۙd=��d��_{
캇�>�:�
��-��0��N�wKA��;0̠� /����X�4~v?g����d+�A�:�\�>Y�uVc,��IzX�&`6�wZ?��i���
6���ҩ~��d��g���f��[�<�L�z�F	�����8i�t��۳����~{]}n�js����z4?���o��T��5�r��Fď���,�@>���&�F�Wն}7� N���m�r�7�TjG�<�g��ɻ;O�R_�ԋ���R���	-�xZ��@Td��&���݆�	��޲��µ0��X�.Lzο�l�mb���L5��q$o/�����\k�AY�~����.��/zr���/�ihn���*��+�7��w��B�@�@�%�W
Į��	�/vA��{R�Ψ�`�K���L��������G���PD�em�x�k,�c��_�䆆����������z��v���j�3rxT�0���4����_+>��`�-.U�T�{7�=^L"��å=f�lQ�U)�T��V��m�S�n�NP"��{���>�<ޜ"K�� Y��_'�e��VЖt�BIɡ�/_c:!A����d=��£���ԹE�1����\�]_�Psr+o�6Ͳ��]��W	����Oi�-8lF�9�Ԅ���7��K�-��v��AEU��)6���M	����}��i���=�m͌c�G��f��\W���)}����q��G/�6��vMU�آ�� �V,A�+K�'�/���;p��{T��@y���4m��do@HTW��;+���/p�N�H�g��u]��E?��[Ϩ��ח���4�N� (����G5�
�r��� ���Z��vz�C��y��*��>d�^�o4KV�����.��M�׾@��gL�����<1������?�-4��pI���.�1�б�z]\���A�bO��� Q-���Ƅ?2���S�b�6|872���ir#��H��;'�b��c�>.,��������i�[)���n�x<�B	�٥SY�h��w�aÈ��� �4����t���:�t��w%17j��Ɲ���<�L���z�W��^�]�iΦ"j�߱)���,����'d��c
�"��Y!���U�dᅵa4+[-���C�I�C���)���i_ �9����0���,%���������*�/���H�*�va��m�ϩ1"��BE%z��<v�-���\�j� 긁����܎��xs\��� �!2�n6\�-���O%+(�D��IM�� D�g�R���6B:7��w��fG�*�5/�C�n7���E�[�[j�}^N�=����D���Q
6ǘ=K͗	��R��g$��2�.�3�k���:�'tԇ`�CM��a�N	�ҕS�fv�����e1l櫖�[}h�{�!��3h�6èp؂D����Zp��/#���ﹱ�<Mv��s�眐�{U�mKν�N����R�m>�_?ehU+����@'���&���qH���ˊs�gmÂ�A��ӏ�f# =�_f��tQ����1�Ԃ38Cv��fu,A(�U�4��� ���j��S�sH#�~k����!�6J��%�{��g�p@��n��R�M��"�mF�{1����~с=2:z5/V��}�6�gn�s�ꮉ��������fٌ���GX۹�+r���WK���U�g��_w�ҙjۼ���:�#f����H�mo� ы����� Zl^[�r��`)7k"i�z:�Z����arte}�V/�|�ȡ�#�Ք�V2g@��ݪy�����͍8s0	�1������ݳ��:�E��{Jha��K���Sbw*4# <�ǃm�F4a���G2��#����J>. ���*8(2'�Ħ\��2��8���}5��Fx�i#���\�&ͬ�:^\X�� ����:��QN�wi�׋���t!!�?J��fJa
��hw�_
9�L#0v��=KN̉Д�~�e8:BؚJ�ڪ�����]c�t���L1J�K)|=��D���f���Z�n�Y�.x���U'���EW��"���1�Y�f��6�׷�!��F�)��Z`� W�H-F���L��-H�x����Ҡ.�h)!ݢ�d�����h=����n'�8o�q���퐖�+�=ٞ�+���a Ԧ����ᶚ0C�<3���4@2��Hq#L|��2���	X%ǰ��bU��h{P�L�QLq�˯l���4����bZ���EGk�cl+T��m��4��w�Pd](��B�.I~��D�nuoȳI��'ad!��ui�iڧ�*9�k�]��)�m{���3�܍���[I}-�/�0��5s���e��Y6���IAY���`�%�1�x�xK�铁��CV逍�QqG���I`Na�N�u{O��V�wքb�2��/�ꆅ]�3_��`�K
ik���I�<��DUhѯ��Y�[�B.��ۡ(��U @A[���Y�Dkuu��l!%T�7	6J2�%ܤ鎀m�?�)y��_�3�-�cMWz��c�V��T�Qj�5�hD�糧��_jJ�J8n1j��ԏ*C������p".}'
4�P"$��x먌��Jg�����S
�d�zzuW�z��t�7_~8�4T��^��Γ=�ȫ�]@����ơ��؟��Ac�����"�H�O$&*Y(��ɮ���@���s�߽���!d��C�̏��ߙ��x���!�Yw1M�_�@S�e�T�S­���M����қn�e?dׄ� �F�hY��	-�tPϺ�	Ll}=��j��Teq&4s�E�v_%�&��$vO)�C�h��I�4�*�u!	J���O\���D�Eˣ��騽���Z{�SA$����I�W�s`.��C~�W�x�� �����ú�S��j3���e��U��;�k��F�M��TR4T�J&����3@L�A�m?�$i!��H�u���mDL9���G�BB�F����4�U���WF.�7G�`ZHž:�L��gr�+/�q0S�EM�ܣ/`���~tEWn]�|���r�7�|��4�&r�u&�"�:�����"x�eҤ�B��ule@{zF��6ؕ�P�0�``�nU׼����5ݲ�j����n;Sk�5�����������-_������c^�Hoy�#VJT��o�!�^t��B����R0�/�r�t#c���\�I��C�T�q>�fA��j���D�g�C�;�ܜ�1��{�]�.8�����RM/��[t����e⋷�=E�� ӥ�wStn�]�J�*�:�~#������&EUB��K��G�^"B���ѡ��<����h9�S� �ZmN�PF�����i�φВ��ݰ�f�	>����.���3�]�MmsuYF���B���cKo��s"��X�����_�2x+��!:�9�I��d�)���C�(�XVK���#\c���]����Ar'TA��{JZ�.�̄+h���FhvL�}���;�q�4��:��~�'_��{�&
D���u=F�q����J�y��`�A���ߑ�K�E�.���#Z����ji)����j��$.D��!�1�z��;�����&A��޻�כ�F�C6P�W�cG��2N��H�W���[���vz����c�3c¹[����&�{X|H�J����'���ʐ�/��}����0/:��U�ò�{i<Ez{0)�]v3\z�k�����"1v|� 1nz����s����U��z�oX>�Ejp>ҥΖJa��=�\;��$�Ҋ�H��P�������G]�-��Z���Կj�>����$��n�N��փ�� 6C{'K.�3��9���?ԓ@N$FZ������q~
l�#7��)"���0���?����/���if����\�Ty����nj𵯫�Ս�d�>IL/�J����l��A��w$���������칚h��/5@/P�r<���9�=��/�q=���0⤠Z<��c@�Y^�����l���9�����=���&�Y��O$:�Z� в,t��F�ؔ<�e����]����_b�V9�>鰵B�5Pf2�����A{%��f��B�AL}R��R�4� C�$���. K��Y���	�;�/oŧ�׆lO��� l%��pmSՄ�ǖ�t��'j{��S`���,7oc�����I?
�r���nL�8M�v��r�`_�)���� �+^���1����Ib+��f�
��^�'��}�yV��C(��q����G�f�V"�da�7���k.MAD��R��������&�bZi��[Ke��X��t��v��L���sLw�,���:��٪����7�*W�:L�Uj��[��H�*ƶٛ�2u���9���5=Q�1�;b�O�z�h*�ɳX]����	�o� z���%Ҝ(��mo�̥&.,Y<9�^�*�+�Q f�&��*֞��w�7!��4k��=�I��:y��5\B�5�zE>��.�����r{�"�b��aN�@��?m2�Oe�|�&���>c-d8��]�F���/{P��+���>��f�'��}��jC�zxı����0�=ߘ�M�M&P��x��ꀝz�Ɖ�$@1(cL������|Jx���$������$������@`����W���!sW{�l��"�7?�!��j��}��
���u�p��B^�`��x�A��[կؽ�'N4��ɣ7�T�&'(Ә�'�r��,yI��B-�x^�+L- k�S $���#]Ʈɓ�h�o�8t�s]��-m���.t� N�e�B<�}�չ�k�]��v��Z^XN����K���&A�YD���tsϨ/�����x��湫�=d���b�ww�*��8s��i�"2ʲ'�gN��]|\��dC���"#t1g�L���>B�
�pDz@�o�C890��{�<:f�l0˟8Q�� �}|��w���u�I�+Q��&7>��T@���EyKeؾ�9TC�[g�V:��_�2�p��<m���x�+�\�?�KM	������:|���;����'zF��H�z�����U����o-\}��}�j�����s��&��!I">c�-�2:�ZM�Z^��2!}F,I���u0i��8����^9B�(�N���t,�@��Ca㗖�Ѯ���sh ��P�48"��y�&9�ܗ+������l5zCph�յx��Mv�r����U,�(˸'O�s��{��'�q�P�S D=l'Tx&���lu"i�&��joc+�=��g@b���7S�,Δ �`�'뗇4'!h}d7����T�3@6~���[����D��K��֋R�9�ԧ3���ю 	�9��B/�Ɩ��bl6���d߲������6������⥯U�g}g�΋mGY&F:�C�ݾ8��|���H����A�LՂb�OQ36%g�
��p���T�L�����媨.~{�LՂ���k�N�:��Ċ��㷺��rQ>�Wߏz7����4[�R�/�ސ\�h27p���&�@��ώ��fnw��$���O{}N�0ò�ε��e2�AT�ǈ%��1��������Ċ��UP�C�G*-(��$X�,
��%Щ�h9W��`��[�G �����K�+��'Izl���ZU��Վ��0��B/hY�Z)W0ؒ�i#��p�r�șK)	�`=+�=�#����+��ħ劚C5�]R  ���WZ��:sУP���h�k��@��g��l��>u��q�|~�����;%ԓ\=p�����=�� q����4\ƤN C,�E�p/b���r�^�A��H�i�T���ա7�� Q%�y�����SӃ���3�`�d�Z�����CwnqTc�۬K��>��:��鲜^�FϪ��
Zf��Hd���|�KT�J��i�%ᶪ	�`h��]��5���Ɨpwd%,��g/��%�]0��K*+��[����=23I� �P�%�P��ؽa3p��혣�dr������.Q����'�x�b����=NἛh�U�x%�&8��y�8<0���H�r���v\N���!b�nuU�c�6/��^{D��b��R)��,f�'�tY-*%v,�1
�fZ$���X/wK���䵢6Q��W�� �&��1�/���0�Ƴ m� �E�����M���U���;��vUp�tĨ��܃D�Znd���>���5��[3�r�yH��Y'���҂^��6�$e.���>_�	M�8�YD�e�7Q���M3�vRC����8���W�i��m�a�\\���d_���5K�4N3#�[T(��$���lU{�m����r���O��ex�cڌ��s~>�nȥ���Y��L���<�C8~E��kWm��>'�e�]�/�ӱ�<��;���J�|H�����#��e������V
~	���*Y���rށ�0.���zv�7j���b��S�^�b�"��v/�5`h�o����]��
�!�	ň��nZ��s��b�w�_r�^Zc�{��$򸨫f"�H���ns`q+�+>_���>�P$f�	�5ו�IU���v�[��o"9� C��츳��}��5/���H��c�Z:��;Nj��3dY����P��� ����q�[�2�7�xr4R{-x4HE� 6O�τN_�����1=�FE���N~ �u��F��ߺ�^^]�-qp�j�|��U��}/�I0#��F�J��Q�W�����<S��%�3�ĠY�⨆9�R��[���"��͇���|�fB��brw��DBQ�k7�
�<�rv��A[�6fϯYYKH�\��pV���[�eG~�fV��nq ��|ݻVa�aD��C4	�%)TU�⒉R�_��{j��}|����+ܵ��Q����|����0r9OW����)r���(���GTЌ�K8`�e�ӹ�N6o�?wǎ�\���}��E(�������t���VC!B�SN{���yA��xw���l�Ĭy�l9Q�p\��{��!A�"#0p�ZQ�LX�I����ą|'əI#,�H���_��k�m���@�.�N��n��U��eVEozn:�r�v#���_&�u�1��i�����u�R�qKT["�=B2��ҷ k���##��Y�{:1ck�8��?����n��F1r����Wi��A)���­����pڌ��>�H���!�z�cb$�k����I��2�� �( o��Ֆ�j?�\��#߄ͯ�y���$^�y��c��c�	�_:)s+�7��hv߮P�B 5�-0J����'�<O �6b�F���s���F/>w��A����FV\bs��x~�0E��?�؝9��Ҧl�\�A�p��`�J��-d";օj����ͩ�&�ׂ�g�boEo�r
�8Ҍ_'�l%�p`�ɒ��dnyȶ��(`�a�t����%W�Vo#�=:֪���>��,� svE@,�=Ë[�z�F����az��
�2|մ>z'�v/uݛv�O��*�{���y5��b����:D�"���h&)Yo��\lg>��ħ^��[�a���8��E���C�ք�#4��(I�ג�N�� ���	����M���Qtzq�mj��/��~���F�wt�5�Si����V�}��r�����0���*v���ǖ���-*W����4 �E����9�f~<>N�¶�gX��U��L�����L���^�~~�]Q��n��� ء<l�&��iY�t��K�|[� �w2qW�h1�����x��_�bH����Գ�<<�l�OxZ]��7��=nU����	E)s���`��[A��Jps��0�"��W�Ζ���}�H�"�=
.��'�,�ͭ��fxE0x0��'#`� �0=/Q���5�U��xTH)�"Ǟ��\|^�pk��]6Z�F�}�^�<;}���_ӣV���T��W|�N+�@��_�<I��v Ď^A�Pw�ܢ�~�9�v0���b��LKy��cb�sd������۶E�зy(z4ج�@����#/�ż�'	�+
&X���d�(���2T��8fZF	�.�ƾ�>��N^O��~�T��k�U~��۴����F%�}r�h�D�X�
Dhu��ss_��Шڹ��D��A�$�ڵ�6�ᱦ$�V*厱�KvK��&���m��.��Z�����/����mwz,��za
��_�(=�\�xl>Aׯ���քe�!���R�*���7�t�~Y���~/��d�%ǻ����B8V�WqZ�p�p�o�fɜ�Q�iW���X�1zY��C�2�c�ɟ!H��O�c�u��ƪ���4y=Xi.�Y�}13N��[7*��/�ɵy����A�:U��s�V��ň�F�Z��| ��J��Kn*��x�SȔ/�3� hn��aά�b3?62+�8R5 H��3y5�_{6i����jW̙�Y��e�e��L�]������C6�Ԏ�3j?����)j���	�q���M�����৮cR�v�o��gB`ė7Q�|����0���/��6��R�U��������c����@)��QzƮ�&�qL��6�Y�KFY�d@�l�M�u+���L0�N��]�	���V�(�MB{]�V�$8$�n�3v,�u����m'��D?�f�ս�AџY��E��BI���#��i��
p����NɝuP5�k!O���}�%`*�TD�F�\݋�0c&� �}l��c`��Ap�D�<x��jg(�M421~�Y"�~�`�*��jDW���
#������ϸ��(PV���,^h�%A�f~U=��s�j$V_�fx��v*8�?;�E�h���}r���Չ)�l�vy�@7\r���]�����	��
/��l�
�4q��F m���W�e�xE<Hv�|�9�-�R�M�J/V>�K/}٧��w`^/�?'�1����_���A�z��m���˚Ș���[s��'k���AP��@�P'�);�2�l���^ysϭ�@y��O6n�ڠEb��,"��3�a%�Lt,7=�q=�u����z�FI�[�um%����u�2�E
���2;΁���(J���J�vLM*�8�����Ry�>]��y��P��;d��2���\�<;rj�R�A�����g��eN�t1Y��"&�@$q�qD��Y�X��,KC
	���j|�"��$w{� �S�����p�ˮ)�ʐ1�w�#���f�o�eW#�:��$�D8C=��I�vy@�hl~d���P-�R�%O�Q�b���%���1�����	E�U�R��^��x�lôQ94`Q�N-����bkv;��)��"�:�K��t4���bm�0����/U�ۧ���������?y~rz�¥�������/�o�Lj�r��v��ՃыBp���!���xn�*���9|�_G�Ư@��yBI�n�ˤ���e4QK<�?e�$Ih\��Z9|*��|t��9R�fv�}��v%�pV��<�md%�V�d�5j�G�G�����Ħ����#*�����lL8/������-����yT�ନ���Xh��5F�c`y*.�Yg�Ә��/�����T�6��A�3�O�ħ`���h�V��w���I��ܮt���pk؛,� �@A���V5��/��V[��6S�JB(8��4!��|
��b��;v�!�*}�˚�٤w�a�X���.��&��Ϡ��Rq�X2���������$����L}"O!6��f��&�}��� [�%��X��^�B�����+�/6]��ߨy��"���݂n<=0fp�f������`Q����@��$�����
�OQF�c	�x4L]:ֽ�Mp٘�`�Nx�]�Zb�\]���p�\{�:��
@5x�����C�W�Ʈj��UϞ>��j���_�'�!Ј	kc��w��e��'6��I�=�G�· �K�R��-����dİ�8��x�X1�B�㊮ͦ�5�143�8g	�6SfS�Z�@����2���l.�}L~����@�˥���s�.���.h�� �~+�w��2���N�e|!~0��t��2눻4� p��\����`�|It�
6�e� -~�ޝ#��7�� _�_���<�D�p��Pƣ�=�&2�x|*�1A�ȿ��	T� F;|j� }�))XU�)��m6�(I�����߭TsLУ��`���i\���{��M�K�c��?�	��w�)B���1,HP���*���Em���ƀhi�c��S��zR�` rr؎oXZA�W�������!��7�q��$ "�}��Hc"�*�E��8��u`�g���0�zŮq"mv�C��X^v��kIp&j4��2b�I�e����v@��5p>i2���V��
S���0�C+��5bq0�H�Ɛ���;��/��[�|"v�>�Y�c��B7חe��*L�G��A%����HdPy�hC��ZF+Y�eX1]�{��*�����)ky��]B3'�|0X,�?e�I���7��ܻ�wg��'���'��[����f��/�vR�`�B����.O^طl-l̯�s��/�0�@����|�P�P���]�BW�)N��ܻ�O?�ߓ�0s�簰�i�?��S�:��J��N����)xnr����7]��u:��FU��2�QzO�ێ/Z/#�j[O�����B"�[}ܔ��̫+��d��#��Y"�_�q�E�;���F&��E<A��W���c��妛IK�U
������v��1D�/+E/�[��l-`U{1����W��Qb�<<\h��r)o�9�.ZwB	�|\�E-�/"���N�E�l�0]:Y�턈����"����j�:qۉ�1�L~���E}�Q̈́������>��9*夁
5L���ϙv_�6���O7E�u����>45l�+�0�D��~#��M<IuVf���X�l�U��2@�������4��r'������5��Ғ7f��Hι�z9���T��ݚI^[ilq	�4Jz.�w����U�N�����p��g�e����	����b�;�p�k��S
�F�u�sC�oD
5bdj�O+��/`#�< A�8��H�!=�ax��M���tUFbj�<'I�'	mh�a
N5Y
�k�Ӎ���!B)&^�Ll�*��n9��
��/}�s��~S(�<}���]���Ȱ���G�T����.j8�P�����c��<R�u�_1KF�Ѯ,��F��CM��l�6�"� �'2�";�an�f��G�V��)Ȍ�9�E)�<�}Ջ�[��� ���d�2�R�������#�@5�|-wtݎ�%:�C��BL��Q��2~%�,��'��M1���c��T��K+�(t!�N[{�m�-��Wɾ��Pk� SIʄ-�FAq��S���:���Gc�&�Pc�g�~�!���SZ��Mc�����1P1]_��[˒��� 0��2-k�,��=��e����M
�l�!|����=��3b3.&2��b�vmy@�{3�	^d��o S�3.�L��B�Ѡ��2Z�S�],�^\�3�����}( ��í&8���T�h�S��;�`/�i����]�W�C��k�6TzRe`��8��������k�Ò ���X�F��[Q-����庅5�O���!	c8J&
MZ��r�}��餠)�^Jr-��fw'�)�j,'�]]���fv/x�tnw�UmP�fݯD1|-r��h��6�O����N��J)]�i#@4�c=��P|�R�������'���]�FL�;|�=����*9L������{e,*��.��o���,���h��w�Η����������U��w~��X�d��EP��+`ohKj�+�gkpG�̜$L򻐱1�\j;.0{�'�Z�Q?�L��na�1�T�)�m/�����`�9DA<����_�Ü`��p^�x`p��g�Ӑ�s�֎�`.��){�h�K����յgӵ����6��Ġ��d�uSgG$vX�=�z���Q U~	���cr�G(���PiO_�8�%3�}��ClஶU��1ݠ`��`�UƱ
_Ǆދ���r�S���ts4�Eyr�c!�n��%>Ԧ�����C�hz �w�-�AO.�c�dr $�Ÿ�NC�{Rȟ#��7�T��\��A���h+����>^��!pr$yX����I[�Z|�϶��YR�.N̬�����Y��EA���P<<&�|����3�B2ި=/Չ���t�+A�c@R9a���9;��q�|���I�	��Mv�U�5�$w�������:�Z�6��2
����������2ABZU�^R��X��A���y�-��a\Z�h�*��-��I�3�3�,	K$�Ϣ��Rg�+��2��->D�k�����ID�p]<�)^S��1�ԘO��~aa���(���@y5QYը��27x7�C�@DT_�f&�ڊ�g_����$��l�+�g!��^��t��c$���B$��Vd�}��PF�"��&�a��'2����p�	�[E����3	�$D�+�1���7�hPK
�`a٪�x���z�%�L�ŵ�8��VV>���Gi��7������$�:|DN3��o��j����Z�\圻_�����[�}��󢕛~��}:w��+I����) �'��=�n�x��?�1g��,1�2�]g�P48����"�LyǊ)��'$R1-"U-�*������H�y ��9n���5�uu�Tئ~��������2��}jd�Z��W)&�ěB[_�ݡ�����F �&*LV�[�C���w�%�ar`��	I��1#�=�OOj���Kً��<$�����7�E��<��#]�֒�*e "��S!}�G*��6;b��4� ��D��Ԧ�tWE�Ru���?�H`������9%T���iEPnepX,��!͌���~�a�Ȗ^�8s��x��O���KtVhؠ����Q����O�}7GU��J��GQ${O��@%�fJ�>�&�b�M�7��,>}����1��ܯ��#0�v�Oy�e0C==j/K(VA�k��� ��_���w�{A��E���l�N�(��;���aI���?�@�Z�5�(<i�IqֵGzZ�#ٟ06d�Ы9%_�4�~�e [����!B�)KABZU(���[���P:���x?r�X��"�8��uX�G����2�(s�~�g��OA-���vs�p�o~�8`�>��N�7���hA����\�P���qgDdե�A$��u +UR�2U�����o�Ibl��;{}F�#����>�A�XT���r�� Y=����?������$E��7�n�2kL�J.�l):���k�R�+�a��Wx��¾�x�d�U���w�m��6�_]��A��Y5b��rx�fʄ���"��g^��Y�/�`	)`Xs���*��욜������;ka�mpH��{�ǆ�V�PɗI��������އ �̲�H�E+��(�%R�&��UdQn ��&ڦ�S��e���@�+Af�d�H��$�z��C�1�&<�����m�&U��N}�"l��;��ĸ׈�'�d�a4ݮ�/��0�D�w�c�ن�	W�q̱�w���A�[k-��	��C��+���;�is�ۧ�Cyݎ(�~ty�~���Z���R�}vQ�9��Bq��.���`��F6�E��o?����v&�%��nT���?MT�<|��B���t����R����v�3c�?���&뽿	������TK����2�)@}�Al=����ii����=�-J-��2�gS��FiT}��\��x����O��k�B��S��:���o⭬\2ٟw�UH���.dt�b����O;���D��_����3��S��E(&mP*JK�v�����_�DE�'!���S����~l~u������;A ����m�6ǣ
�=�r�Z��M����j~�1R���!&�n���O���QT�'�^�Hyӭ���G�CI�͒u������=k-
�T�f�$�V�'�p�-���x�g����b?oV)ؓ'wF�ea��^��p����>I[����<
���Ķvo�:5���i�e�)��=ƿ�4�3;���<fk��N΍�0A�N���f�Db�n��V�λ�s� L��B���?�e�g�R)��hVv����KbG�(�����(�J��Hov�����u��Y������+�	���q�?��ބ#nH�L�o�xJQ��}����#a���`�ĈYK% ���̓Uy�[��n��#��eE̍{��(�OA��+RS8���q��̆�N�;$J�߈c�����>9<'Ս�v�8V!�p�rm�f��>�v*)�tjd)�͛� �P��O�7w���~u�21,����=Ĵ]2Iƽc���{��&Ղ�F"ŉrZG�vr�R	C�k*UP�yhpB[�C�	ev����������SWsF)"����_?��eH��L��X�+j��٤Y24�?��z�;�v"��a}jZ�P��Fd]:�ٜ	�O��W�ͣ��s�Z�m�N8�LK�z"E(�t�O���#p����>��4��G�@C	���Rx��d�F9m�ؿ>�ma�RŲQ4�k�>�
���Ӏ�r��[���"��D�iA���/n������R,%��7�����E=>��B�C�	�hs�\|��Zz� q��x��!��4.3t^����o�=�j:�w�\=�?К(l���R924��n���`'|_;Q��j]�}�v�����P��D^���ȝ�_��,[���+f���nZ���~�2!�#HƟ�`� ]�S����v�E�s�ҡ������e�jnkA��n'���n(]�o�R%,��u�l#��}U������l���Z>�����:g��t[1�F��/WWɷ�h�����j����0��"��fȃ�Du8�׉�u2���C���1Mls���Z���
�q�rl�X>T=Ve9�@ ^.m�/*gwήpſ0��cXE�C��c��FK�%�<�$k���)n�Xsd�Lߜ:��8>nF��59�1��+���UW��J����579�W�a&ھ}#��@��߱�s��͛U GT�����=�{�b����@}�8h�J��{�C!�u�1�~"�"���>;\{�*�ƪ��@���:|��,��s���7�v:/2�?gJ)%���kLj�/�
���r�<�P�"^�n'԰�X��&����в�*$��A�����v���~mq?������cWLA���ESw���:E�Kv��
����Q�J��W2�.�*����ߕ{�H���A|	��E�;a))VTdgb/
����m yOз��͇��{I,�1��ɳ=ԩ0��U�+D��i����k�/;.��p _\�<M� ��[ 
��7&V�T�%CS1+;�H�&.�5�%u8˻S�zh~�:�pH)�Ei�ˈ�g!�)� �S񫏦�C�A��C^У���Ik�#:�����Ӓ�ll~�Nx0�0c���}�0����βaRgg���-=k�G�辨Z�^VQh��e�`��$�*PGs�
U&�$��|����9�y�lɣ���wg~o�����U������4�nH�WA��Wl�Q�2����w���-��5ː��5����e�/<��:݈M�]�c6��I��`vn�6�?
qx��[�5n׋��/c`�kݦ���^x���'�x���)4��&�����p�lȴn�-V�Ak@	�n)0&�O���#��.vXĶ�)˻;ִ�i�U(�&��L����d��-�}`+[	?����r��;?I�:��x�(�m0��U�)��7�z���~p�q�눎Je!�~h�K/wm˥��U-謤�%̰gf�$2���hA��n��8R���<ӵ~���g�t����6e���~ �һ ����7��1���H��ID�h�*�I͕��` �Q��I��=!�J6�Z��d�x�M@��|��X.%㚆�p�g�KݙB|��>��4s�:o��L\�f�����^����4@e��1p�g��J=^6����*-8�tW���i�qQ(��s*:v� ��߱���]YD�٤雁Z\L
:�#7��7ɇ&-6J�'*���Jd�L:��O�$�t��F]њ����*�>�@�jx�oѝUs�~�^��^�C�Ə|�f]:\�+��֓��Uu��N���W��?ac�"v��#�r�vx���ذv[�r:`)F0ܧ�g�n���i����hT���S�̬�r ���įF�,�G&I��tt�z�ŶRn��S��i8�GE�(eǓ�hɒ��R\U"鄬��U���9V��6�/�6|e�6 �?t�H���O.���_�e,�Dբd�8I�h�D��f `y6���(�?�z��U�:Y0N?A��aM�[�;�9�C���tl^5ʁ5�"�*m9�Fh*,�'i� �i�}�����cp2�i~��S����w�5�,u��a�"�Z�5��**�㺵���2�9��BGVa�I�pz��9̏(,�M�p��`��-��5�CS��n�\��J��5V$<j���q�P>y�.���7y�йآ�!�,9|��8ed�h�c���!��P�S��@h�XT�8|c�є}5?>5��Ow
+
K�U.?4� �Թ�:r���^�5*
�a�DjAu�7,�����A;h-Y�3#�V���)Y�0e;7�ʜ�#;G�Y��F/cl�>ݖL�6nAS(�����JsO8�*�<v=hc�^q.@k.�Ps#ޅzU��ӎ��rya�!#cms`T�Φ�s=���'>cAYm
��m����#���Ry)���k����iE�Ł�Ӕr�?��_u)�}��Ƽ��)�{Ӽ�q ����P�����vo����}�zֆ�h�:#l���!��W<��. D�lB�I���ZSD>�Y�V����$�J���u���g�堈���A���{U�z�g���sȋu�b��G�E������091����6�c0�c�'�p���-j���V6G.�9�K�]�T�(�G��>�r�v(������m;�W����P?[�k#`:����A#����z�e��e�Ȗ�y-m���~�K��x�h 딆�h�_��h:�^w8;$�)j�C��N�q�G�yPM��.!T<�M�t(9�O�spI�-"\�Lx�����Yk�l�o�l�c��� �4Fw߈�2C�]�Z�j��)�̫ȴ�{�B��q=Qq7Ŧ�RL�;�(o��&7bxe����a�t?IdH�{�7�����������q'��:@��?�ݰ��C�R�Z��6'����I��˯X�5u0�,��amy��9�����E4����$ � �DӲb`�U�ī�!��٦����'���c�,]�l���KϞ8�,����.�x�9�HWzO�
��#�N�9V\�	v�7}bv���I�,�N��w+M�Ÿ�kp&&��s������Қ�D�Y@�
_�N#*��"*?��'~�����jsA�YN�ݒ���x�Hs�8�F��eC�ڔ�$5y��am�q�`��Y�
Hp��j�M���;]�a�:�*T�p�M=Ǽumf�z����Z�e�|���Z���	��Ԋ����C�7�2\�Ѵ|�:�g�ܚ�gX� ���ĺ�%-�E�6��l��Rnڜ�xU�Qr�^��Y�|[wB@ʬ\NNG���������d���v�7��9>��RYh�ͩO�V�.��#�ӱ���&PUl$����Jp���
+��R�e�9���篓�s�fI~��ؒYm��i���r:�����{�"}��n_�^�k���n����+����B��ЫýOh�4�f�֓�۝)��Ze؁�R5Z-?I!�Vk�t��m�I:�I�_:�!QJ����D�"@�3,C.M��W�"4}UA���׏��Ϋ�$`S�׻����ߺo�����<������nl'a�(v�߂ʦ���c��d>���$�MW��d�����h��4�fOq	�-�c��F �l�B���O e�bis�x���)���%"a0�
FX�5m?n�	�y~;E�_�Lr�,�^o"2�}�Y��[��h{"�����>K�Ԛ�.�%�a���f��YnN��r%o/��8�!��_�Ag�@�zyX-��0%�>����V&s�p���<3�Y�5 �A|Þq?�z��jW$%����8���n�OH1��K��&��ӿ��G/�/neI@�A�ə���0��0/�͡q�U��q.p�6Hux�GۏɌ���,�_�C��Ť�˪�q��2����y�m��A���9YGߕ�n������A(*�PAyr��lvr�{�;ݤx�-B��3��|�cA��^���|g����*VrS\�0b���\tsނ+��<���,��c����o���C�-U	��Й?�s���L���k����ڋ�.*$�z�7d�rƿ�5ᕃ^����O^e��x������[=2q;$-�ք"�ģ�Kx+2�����h��:��W=װ�5�sWK��t����&M��HSk�N�5LBD�]uo���Ż�B��8��c,�1x7���}�J�� c�SO��\��K�*{z�C��Rz��������XNb�i��,UW{�p�ic���msM�T�L?��8�[)�����"�v�"�r��n()o7��@+�_��矋
.fɆ��E�@���}����#\,�N���{S��[�j�ΒI�i�x�5 ZtK��;-��9t�C����un�i���%k�������
�|2�y��<�3"#==V���~4�M�{J k0�����F6=@@������A��?}x��]�wp,-��_��q�ߛ��	O4VmI�����Ȍ{�HD������ͷ:דꆼ���X���pRd,f���&��Pؓ,�<�w]<9�"X�G�+�½�R� 
|���,b�$��O�R��%����
/���}O;:_��Ψ��,q�P��@��+�;7���gFy	m��9�|�0��3���z|1l<ܙP�S������jY=5�wֵ�6/�����H#�0��'�;H����<��j�0U�=x��RL����(�T�+j.��x�ޞW���&�z�����z����%8;�m9�,�ښ�8�o���Q�S(���)�؃ Ӣ�\�ԿsQ�sg~�h��Z�y��D�[qU�`Ҧ�\9��e�m�;�rN�0Bqٌ�D*�yv�5����j�񒝥6O�18���M���S<���oZ�[���e���5z�����>#��59=�-���
u����ĸGQL�e*f�6a�G띬QK�9���f�6Z%x<�S�x%�g�~OW�4E��W���r��-O���y��/�/5�F�&����nQt�m�����@WM*#�����fBW�Kv�H��.ib�q����W��R�2��)m�hDsQ�Y���d�����%!�+Cg�D��I�Vx�s�B����.st��^�����\	{X=�cW��z(���7*/Ώ�W2��c�w�w��4��������Y8Q��h�	ډ��"d�� ���!ylaS��r�d���T(��{JV���0#p:� �����/n������&��IX�'�ȳT�4p=ͭ#նtZ'���9ѯ^�<0�+�4�+޼���V֎�����F{bN���_��5����,g�Ĉe��9�k�9@E~
��7|�n�9kj� 3U�	 �ohot��9�*4m3�!V}�<�ߑ�rp�C� �^r<��U���l���d���)
A��\WF��a �tO��At ����@�� j�]�k?�x3Fq�'#C���ĸH�}���(Qdz�x�$�K�W%�]a�hԑHJ���m��b���qC�7����q\��$�#ܒ�����.h�u-#MS4�^ �Saɫ���`���>;ۥ���);e�1�Ώ��T]�\uZ�Z��*�j\�:E�J���f��q�E�V3�XC&d�	,��"ʪ.*Ƥ[���ϭ�g��׍��2-�Ǎ�c��D6�+ �u�Hg����cg1�s$��� ���jW��%�e�t>��n܅�j�CLomP���
���M�p�1�+�-꼯���I�R!ߑ�V�su�$����
y�O�������*�#C�?��`C��7�Q��#ib�k��<\����-��>�捴"4�;�Q�ˇ�C��uۙvI�q���F��$�`W$t���G=&B�B%���%�I���m�ȃ����g.��oq�$m �b�H���"l6>��@*ϯ���@&���s�;Y')Uj8�+�9A+�8z��䮒�A��C+�B����g!je�}��s}��^"f�R/����1�#�kY���HN��`.�0�c��3���+��n�!��ޮ]K~�>�����7!�R&���I4$��t��OG��P�=ƴ�M,J����n̎�U���u'	Gפʹ�N�]Oh*
\
�1oC8`S���nX��0�qLN� �@�a���<�گ�_��|�0`�N�ȠJ\w����E��Bh��2h�P��􀔟c��()�/�H7�R��$l�L�?���%��t�8�� b�;�ͬn8��֐��G&H��+C��ܝ���^��y{ኽ��N'���$r�5S�)�uT�6%u�q��R>CUg�7���W1Z���Xg�K�߄(h\��Vh�#�cT��m|pQ��c�'K��7�BjK�h�����A2�ύj��rN�9�&(�vH}�M�̋V������t��:�PE�gls���ρ��?Z}J��Y?g�Kt8��s���ÖsÂ����U��P�B;�X[=A��@5�����L�;�$�'���Brx���� ��1��U-���vRu�3;��(�)��b�>���i�@-"�(llv��}�e{����xJ^ ��[�|5�ȤwWZ�ִ�`������9��8.�M��<����vZ��PkK�����h��=�;����W���d?ZX'q���#pk��l�h�����-B�-&��@ƽ�l|JW�N��	��nR�A֮xĝ�@�`k7� ��|4���q�����'�sB+�:�-Om��Q=��hT��OM��>5����_�*({�3$�.#(n� ?�becZ�<	����?��<��L&� ����c&��y:87�CWx��c�'J��j��&�Y��}
3�s�3�%+N��im�qf�R~��v����)\�F�%���${h�������!��f�!��@!�N.O4��W�h��Q�R���p��c�E:?��QT�&U9��2@����v���T��O�n9�7F	Z��;�X�Y(L�j��k0���v6���V���˥4��++�NŻ��H|z���h�8$�Uֺ�v�U{?�:3�n��ЌH�U��_�n �c18�?�o����6w�������f|n���ۍ@�00^!�#rN: ������|13G��Ē�c�4T.Z���\�4�g���
��Ts���_ϧQ�$���|贖T�8P5t����\��%��f
�P�����rs�|��s�� p�$�rVw���TmF���ź;��?��v_G�=�Ҷ�����Q�z�x���2�.�th>�����žY�r��
��t�@ �}߰�^���D��2�4��ੳ]���)����� y+��Q�U\�o�9�����2% f� �lЋA�h5a��N�Уr��:J��CN�Q���5Y@��au�D\����$ �=���5B�N��ED� 	��1=O?[���k ���9�*�xG�V$?�Yo�� ��5����h�na��g��jl�;��O�����T�5��P�>D�7T������$�bÃ��+K����F���/�G��4���ͳζ�ж��n�9��-kݕ���/ȴ������_/6V)$l�Tz;N�d|��I��}BF��
�:���B9G�Q�Vt��_8������<9�9@"p}��"���
�ݹV�串�G���,��V>V��m�dNc�[��(�d�8��D)2��*`<t"pV<Z�SwS� ���R]�\��~�W�~��Y-?�%� ��-0?pQ�>��^윙�Ƽ�P�mnHTha��+��a] ���#j0<�Ra�j���ɒ��qٜi_�@Ip�Ԟ­� Hd��X	��IU2�S����0R��T�ȼ�hO�������1�<+i���,��y�g�7�*=︝>[θK�& �=����ˉ,�A�,4SQ��.H5b��Z&�&u�j��u�8�K�h�t篺����n��Y$����Me�>�1O�T?�S���޿N�CjG?ӫ,�@+=��^�7��������3('N�T�z�?\DS�D��7(6$��$��h��5F���T5p�{�464�\��qm`ȥ�8�n��j?2��s����c�,��7p���#a5���@V�q_�R�@�a+��5=$�ũ�@vI������.a�&R�;Q�h۫��]����O���+'��דԮ��{�|�|`����B.�a�m* �pv�)"$�^3��g����]׫�w�Z�9F�Z��ަ �4��PMOxI���k<	1���=ꋑ�CRЪ�1�d��)%����׃��T�8��?�h�5�j��Us1�xu(]d�����%�CA��4��'+�{�h���1{�;]&d��,�0F��Z��k[>@$�9���!�!h��0�F#�"D��3�XD���e���P�SL�}W��@{�^�[��VZ8����I���b15-^op4�V$����Իo9^[��ڎ�	ҼKĦ_.T����K�i<��ɮO<Rr�l�J?�W��X��z�(��.XF":����!As����
W����iU�/�g�՜O`����t�3K�2�B{�Xv�.M^�,��z��W���MC�>%/���ͱ(Wt�1B�8N�9�T �	��4�.�n��	(����d:�/	�B���JM2t�M?�{+�%a�����$��
3�'�4C�o�t��_#=ؼi�ź@SGrk��� �oc�
�������D(��2���b�O�OVP�^�>"|Oi�68�w��>��̔�&���{H���{�_ă�*]�kW�Pj���k_�%�*J.!S�ɇn�ַQ8AY<��~0��G�ķ�[l�D榤��;=@�V��#RC6��&Ϡ\����!LN��&^q+�����7_��Op���YH����`����;�w�d���p����u���eb��(1Db��NZ½�[2��Z�v�e
�l��T�|�M3@lα<��aʢFL���ox:�|���E�=2�ȕ��S�o��6p4�v���N��yj\�X6��l�1�/\j�\K�J~�f��L���,&GZjݤ�x��EOT	y,.?i�w�\V�j�nv���PO�PD'8�4y�hyMN��핀��+Ǘxʾ���-�G�e<�w���XI�Xo������E%m�����51�><g�Ó>`�+.�1��Q:L�����ڣX\������an`K��:^p9޶k[��U}r]����(��������E��Il�t|�_fP�Ƽ�$���!��F��'7;��T9�"�L\�Z�W$Ʃ�+��;q$���QjyE4ɻ�jV<�D�����a<��μ*���A�͕�fJ6�mQ��̏QS��<�ʧ�>��w/�殖1MY4X0��~��d����]l^
�`1�N� \p����L�M�x�r�`-jU�ƞ�R��.��J�b�H
��w�Oªs�O/<�����xu	�x��E�Fx$�*/0
�3�������>�?����'/9���ɉ������+Fbjr�@/�Ai"��0b����8���HZc�8��X���N�����.����U��� �F��`!��̞��X��%,��b�[�;�{�F������ۦs�~����?Y����M�Gs�-��^m�"�[�>g���|QK��'�%�F4A��sɃ���M�Ș흈h�	7�]�s�e�i����D����:�~�
�kX��{�\���1�Jz؁��f��*y(���.|LA�ͯP��A��Jj���A�3;����۷|��iY�az^Þ�����j�Oಊ�]�<YH�}�ǌ1rf�8Չ��kO��g��s�e���	���䫍��(M ��	���0g�����.���5�5r :p�S�̟d]�%����/�D�R��u����v�ҕ�Z�, ��1:��lhyӼ�y[XG��L�`}�w���(yn!i<+��W���㪳����WYv,x��G���.������Fs����{~	O��c�V��)�����ԃ�Ǫk]k��hOG�x�Y<@>-�L�+0��;��Q�
q.�8�s}/R��B\$F�m��Y:40SӪ��n0F<�?t �0j�y{�}`S' !;�PnB��E-�t*���{���h<3�<���2�,�M��s�\y+Ƶ�3v�tzE�� �e��H�m��@�~�����K&u�Q��.��k�E��A-�ll���#���-�!���Oh�J�r[!��ۆ�����};��B�؂0�8O���&�͏
�\\ϑ��/P��.��^�����C� (���=pu�fM�r�tnm�=�Ǯ��W��Y�ۈbi<��5-������rZoMoSf�4�T2m��d��bH�zV����f�m���i#r>C�������?]��p���-��&sN�6�I�X�?��r3�M��㘚��ϖ���,@�{��Ik��P eG�#�2��قU���^h�.��/
���L��k����caC+
�6�����w3�|�����u��z�����kR�hDMƋ�
⠑%�m�0}���W����1L���J*�r�?���~�����C.�TaD"�t�g�Y���t���W�[T�
�+��FK��ҔR�9��T�;Q���|4�_��zM�a�G ��x(dΉ=��w�j ��C��G#ppǓ)1"���>�43Y($���Yo�~9�L�S�׺\]5��ht�M����g_�=��i�ǡ���za2MusK�\-52�U%
�K-Em�(6r$���H�z+~��~N�w�M�C�j�6�K�HJ��`Y�ɡ�+��p�(۪�)�6�r�&N��OW_���Il����RdG,C�,2wMc݈�DKiS��1J�!률�:�,�_x��f���ZE���=${H�.iEXԃ@O̧8q���q��
c�:4ԫџ�i ����.�+P�ۉD����%
d��^����`�I��>���?+�Q�Ӱ9~���vi�x��4Z&9PN0����`�o���d�N��l:�-P}D�`ة�+��q���Qx|�J# �t�Z6[�1'��a?U7�-�Ǳ�����|��c�<n��W��"�̪U���#�R!-�k���1����#����]7c�í��+ނ7�jI�l����� ��O�e��ُ��zAn,B��/����Kg�O%�$�Y 0�4Ӥ�r�El(�^.g�[u���C�s)J]�Y-y#��|JT�?��-�牯����10��.���f�0}�l9�}zS�8&�?�fDn�i���2����'��]4����	8���Ʌ�4��Q��f�� l�<����l�O�#?��Y?��[�����e�u��4��za��{����x��)`��^��m/4pA�"�XAr�&H4����z�]s���L�� z(�����J�������Fau�H#�0���D#�d�{w
@�`��r�TZ.��l��k��]��
��?�j�l����Tuh'w��2xb@1��d���9AGĚ��>�=��Ԏ£CO��}����T��]��kK'C݆�a+��
ϚP��7*��x�C��&w�"_���`�������f#�L�$-��n#���}4YbJ����d���GNE��Ea��둛���%F�,��s����15;;	�F�x9G�@��Lo/(��0 (�5�D�g��@�?�h�I҈��ʇd%|��Ea:�
6z�������t����-:��Y@(CZ�
�Л�Y�����EI$�E�|z"ψÁ�����8{�;㟭qyb��PRm]{4���B�T�S��)��_�>��9�>�j�O$�kD��W��AB�j�r������J6P�$� ;�:�e�:f�(���0�0��fQ"i4/!�^�bOw�3}��>�n@�-{���y6�{���R��fc�VG�zOn&	�ҧ�~ L��/��6
�y�22	P&#\�ü2�zp�����K%����%˧�����f�k	��b�������x��m�QJ��ސf����`u:r@v��ieW5=��isF�cj�&����N�4$�e,6(|Y��"S��D�(E�&��SWp����A`����s���	�ɘ���E�QQq��&NE^��N/�ѽ溶T*�s�ҫ��{Ӧf��'�y.�qL�A�:�65��xyʑU�BN�Q��wA޹�_2����lp�1�)�{�����fi1pн�}=?R�)PA`���~�e�;������x$ �k%����]�t�+�#s�����a�N�7���у�5���ȷ	 �3p�|#� �M^W�M%Pdԏ)W���"GfƜOw�p�51�3sf�/9e�-������9_q8!���[��@�Jʶ�@��q��r �B�3�>iptD07��R3������A�����,Ι��:ϳЌ.�� fknb�у���h9{o<#�*2�6^�t%|��[�,�"��S��:	A��	v؅UPis4Y\�RF��X�R>d�O��ňd���C�dkT�� �!I%�tph�|A���Ծ�4���󰊴׷j v�3r�s6U�t*8��F��ٯ�}��
��S�;�]g0�!�ݦ�O��c��x�b��=�S�^h�nW�U`��p��	������tڣ鋁��� ��\ K�wK�?8ʗ�ڸ,�ȣ�v��p�=�"�L������â�����G�`��]��ƹ�.��܊i�������X՘�+�;]�Bk�z]vȍ[� �zyV�"G�d���D�R��3.d��E�j��Zg�<���X�e��>�=�E�[��p�I��*�-�Z�A&s�J`��P0ǍOǸ���N��x_yXǋ1�lȼ΋Ǒ�N���@����ONd*�c��O7��qԩOᘈ�9 �ڷ��^���D�����g��|���V�0հ6���(Jn����}����m&#[  iK;�<��f��I��"`���]<�X~����gcr�7JX�^��!AiT�	�:+��K�+~����U��C�q��x�DFf?�k��]���!\ZK��&/L="����W���4E��:� W>�3{�N&�o ���W�E2������6�/0��r�;Ul��ٗ�1�h���W8�k|��{��ą�c0b*o�|8���	_X��J��3��Y ^Y��&W~N&�]
�#տ۰�F#|�� .�{�up9��C������,��Y���>t�+h�&g�����"����*VZ
V �R~�)�H�MdyP2�����$VK�c�=�E������@̳�,FHӶ$\�d�F��3,ץI�"/�ޞ4�n��{1v1��X*�o$ e�8t\晇_�D	Bm���,�=�K)�;eN��i��*v�*|M���`1lL�u�w��V{�:�k� ��i3Lg�����)��[��Źa��6�H�j3��R��a�XJ`ŀ��9�/G>�
۸����NCN���2_�S�$6��m��~78'2V�������Xcu�W�	:�:��G+I':�����3E3;��N�[b��c("�b�M��ꔡ�{4�E>}�
�Q���LV�Ob�������d9����>v�_���a��v�ʦެ����C�{���m���W���QV����u��@:C%
+�����j��>D3�09�s#2n���X=���H�qZ���#��5 _�%GyA1���y/gt���F�'F0-[�0�j:�t��� g�$�^g�<�s)�ɖu�r�'�?p�U��dk.$�ݽ�$�<
�	Ļ��{E�K=����Ɗ����h�\��U�"_�b�/ɭ�5�"��n��S~��U]t}A��ά݈>��Ӡ�$����2 ��d�gV�+TVxQ�?\��)K�*��%4���8��h�� $�q�7bg'j���ȫ-^?�A����G�<��K.ի��¢t��_�,Ͳ�
��6��I(U\Ls��5�W53�D��W��K��ܣܣ��)φ���.�T.����[o	k�\eX�i�n����Q��\x�zLh�jg}'Rc>ބx<*�(�T`����,�C������]�0�9:�!Oʣ]�55@�-V��o�Gj�Ǧ~芕�9�\s����T#��D\�K�sT�$����p���a#�p2)�v��5�\���@$����#��a�j��t�u0��<�4h��<:s��U��A�ad{[Q�e0�G��(�H%�DG�R|�]��4�����Ta]��T#��t��)"��";�6�4�g���%@�[���Oa7�I@&���d}\�8Js�È��%��j�N<��M���M�xAj�/�tl�*{�V�l/�G}��B}z֎ϳF��h�eJ��c
nS��o�΢hd�$�(ײ��j5m����ӻW������&�*'(���^!tȑ��� ��&L��f��bK7]��P{�N���E�Au��W[�a���2�]�hkh�:��3�?�7�k�5�_���Z]�E�<���e]P��g��56�H{�l˒����i)QU���\��:��)�	I`�ʣ���� ����Fa���P�`G�Ο-�S�h_���`*��5�J	�X�o(��{i��(��� SLM|l�T�T�!��Ӊ��Y_�G-�ɹr��z].���cQo2v���,ƹ���}��?hz��2&ro��l����N���M{�O��q��hQrG�ެ��P���~}�����J�;�x؊���/����&�HDS@ס���S���0+e�%u��^��H�c�^Ҋ69ExT��lI��O��A�ȕKڞ-8�r����u��9{��+�O��6e$2������cY�X�B]��Y�c�wX١�|�rvMn�gq�����X �
9��Ӂ��7��F�j�=P����3^:��E@%x������-1�������ꏊ�"��,(@7�Ў��Uc��0�V�7S0E����/Ĝ��x�$d�t�xj=��0,��O�R]��Ho�!6Q'�d�L&Ҷ��a��]/�(P�O3�Y�Eqmn��_"������k��/^5te9�O���r��]+@����w�#���ѕK�����[�[�3����߀}��QR���c��+Eh�V���!��,A�'G�.V�8L��� ca��G�pɪ��؀IW;��=�k��6Ը���<y�@�}?�<h3�zp�j�۔�˯��sʂ���8�u/�Is��X�A	�Mڑ��d�7���`C_�Th��DeW�΀�88�%�gzYP	P��'�HfԶ�Ώ�T�@�<�,le^�G�������?������#3���SW�xL.!�a�b �&A�ġf����I�9�E�H�;��}<��,��D��+y�>H��֖��o��U�"���a��l2Ymϧ�]H�:_xrn3�"� ��@cQD%Qh��&�� �����v}��j�D���	��:��`�U(vv̚�z`��0�[.xM1l��4t\p{9ٓR*���s�7�2~���b�D �}��lF�Y�m�*Vh)���ˌnN�����q"��Sc>H���v`��O��O��|,��0G8�3i��")kyP�j����+�E�я�r204�E<1]��<�`���C��k+"e	5��vb���t���[���UKj�B8�M~u�g�%�K�a��$�����VsN�̇<T���v��h}����f����C���3N]+(��nXiׂ-fNO`nH6�T�)����SN�|q������t2�7.�d��m�&2*�S�v���M}�͙I�<*ϴ��&�<�f�,qao�Cz��EL7�����:ٞ!��ЖDN��<��5�/�9;"X�ql�b�yq�f�.Z��%��FGţ��lP�q3� �d"Z��#g��<����³���@�d�.���/��䭐�ȹp��UNq��2��m� �#P�������y�#N��f��(��Bȝ���
ɏ �J��Re��#�N�b���#5��`x�����T� ~������m(�p��u�`�L��NE� p�>��^)$]o�� �y�.��]\�߀ouIYA�D�qn�s]���(n�q�Q7:GO�e�9��o''����������B�D��'�����g�2����9 L ��</D^�IP�\oR�L��?%;���N��V/�iJ�3�doMd-�j��P2��2Ɵ�A�'��e�����d� h/�8���89i��I�i���8��O=����Wuƶ�q6��=������6���,7����Z�Dv8���9@�����:G������P4��������5���R��q"Wwf���P5��˧v
�P��g�w��γֳl?|9dá��6v���a��.��=?��'_�Ͱʁ��F�cC�-6of�ΌGP�q�Z<@���6�J;��h�~�[�Ь��@<.��7w�(�٧���A,�$�`�!����4�P��F�y]�T�խc�{o���5�[�U,U0'�0'���m�^�?��1U9&u��s����'�/�(�^���)���*GoG��@�[����t�R���pV�e.�O��Z��8�Qt� �)������UU=Qr�t���f72��$?�\��?�X�8�"��~p��wuo��z�)7'=WQ�-��flv�?�0rEBuv���u�(�ߍ��8�W���3!�5��1�kC�ޢ�PZU��1C�J�4���pjl}�98�Yn��69���Yt�۷�����!]	�ݓ�{�9�L&H��g���SQyZ�����0�d���9i|v;��}��FV*�?w��ѹ��
12-��K����ȉ3�n-�ۘ�Ș���`ͭ��i����no̴�>�[2�G��휿�b���1P��F�k�ޙ'������ #����@9���;߯,x��~�/ce��|Y�) �$sd��N]�n�����JsD��ԌH�8!��*��$ݒ,�<�Z&u1sWU�3|�s:��E����=U�b��oz-E� ��|�vNƼw�t�v��������e�w��~���rȷ�'��u��H2�YGt�7�:��4�'�{�c'T�s�~SW`n0X�����?���h�`��>�ͽCz�dD�%��>����rʦ�3���~5h	�����_��p�m��Ǹ�vS4�&9���-���I�N�F��MnH9�Py^b~Iqic]���y�\��C��i7��� D�A�j:(�:f�*F 2!QՇ��|�/c�pZ�0u����E�:WIl���d��P4����{�dD�(��r�����]�W޺����gP��#�>x}��!UDDXp��
j��!�6��!B��
8�jt���p�D�O����"�n���*]�=���Q�������ǹ.��U@�z����b>�Y�Y�j�|z�he�g�������\��������=�!��t���w�k�v$�si��`.}h-��# ��`�F��I^�3L@79k��Zz��O�C��0�)f�+�{�dQ�c:sM���%�V��f�?����9	uM�'0�@�<�0�ہ�7�7�_�(m�J�Qʋ�q�����5a,Ȼ�_^15��fL����+�gNyy�����CɒQ3���KIJ�Dc>Hӌ������S����h�٥f^_�jɇ4}��N%�07�	O����<y{텒샖���+7��=4C1Z��mC8�<���b�}:����ʱ�ͅ/&�_\b��u4�7����y�0�����'�a�������%L��>�JM=�_�->��͖ԟ,D�����ws�m�� �)��ߴnd���
o�!����#�N�*x{���V���-��8x�
o^@�[��Tj:�&VX
"��;j��-K@~��]�R�F�������Ce �q�Zp�J�K% j
�
מ��=������ү�:�C�2�M��N����(�쀴F$ ����E��"�k�i�t�U�y(�
�E�P��.*n�)I1
�dJ
��"Z�1�|FIX���ݠ��|EW sw7����g�!��E�U�R��|%�tL�	3a�3 �C�Ϋ[�Gr���|��̋5xp:XJ�m���
��LC�W����N�����	���JبS��Iž�}����Z��)�!q�����`\F-�?�c�'�/e�����0���-戮ÒW/���P<?�p���b��;K��fw8�A��8���hg�m�E7�����d��gΗ|r㘣��!Ĕ�[jT�6��q��X M���.f|����eXNz�x��9ÒO8rU�Kj%v'����Ru5�]���e�����o��3�_KU��о�g��wG�*�Nd�7 !2`;>\\C$
]�W�Ao_f�Ӥ�F��c}3uk��!�1_����/�r�����t,�kL)�ڔ���^�q�C(eRHN7��G�6�n�O-�j q��J
҉����ػ�eUjE��#����4�W��[ʷ
w�3�vY`��)�g�ё�Q��w妷s-�#���`9���}G��[)�Z�l88Sx�X'�AF���}e'������k��|c[=��V��������B�U�x�����{��Uk�:	������n�A5h�b�[9�Bj�~�֮W��U��l�z��/P�	8MLwy�����<�@șҜ0G���t�%��+O/xS$�`�g~�7Zn&��{�����QgIē8dU�\L��!lbW��X%���P���'%+����p̜"x�ԥ��ھ�R�-h�@"�_YV�Ƣ����l��Za���|n���hcl-� 4z͞V	B���k�q*\�%"[�{`W�&ԌЦN�)o�ɻv��d���X	�wOL��V���)��6�?��'����u��u�Lܤ�ԏ�#S�f�1��wO���1��(������\ ��j �j��̄��C<^���`ⁱ5��H��UN��@�I���WF������Τ���w~Pu�� ��>%<������(�y�������L㉻,�7�2�9�Z�b�eQ�h�,S9��-%B�e�j�mL��ۘ�u��e����+4�[��m�������ݰ56�tIF��51ކ0v��?w)3Z	��y�J.�Lh���+r���BT�  j�"�7�gz�K���j�FK�8)\���^��*i{�yȖ�ʹ���5���8�G#����.���&��6*δ`Q/80�y��n#6K��n��kan�Z��tsG���\�b������}��o�R1�_���� �]�Q���s���D����\��M �������� �����~83�!��E:_S�j{0�*� ��t3T���aL���M���(������HL�����z;)�>T�T�'��N�M1��潽�A�m�rfݫ�t.X|ޛ�/t��9��tWI,�2�2{Urd��~�[��z�o>o���&t"��?�X�r���e����gIn����KОC��֘p�m}ǒ���2M�E�u�$����O-l|��	��� �����Y�
Aކe� H]��p���8�{�(豰�[b��RL4��j��M�V*��.�(�=|%I�MO���]�IgԞ���r=�	,����/$���'�LI<Z	n�<$b��e�m�$�9p)��D$�4�3/�09��g��*Ig<3���u�]]T��F}�Faf��?[qm���ܬ沒@�KuI��v�;��C�/.�*Q���jB��X|	6���6�;9ߔ������pp���	�2�埩C�R0�<L �Ex�ds�"e7B76�z�2TV�����i�ɟe�&�Q�vm�̅0��~�~oR ����>ڞ��ka�k��K���s'�����9��������=���}Hn1��V�漤��9�.���g@e���B�����fD���'Yw=��o&��5�qoRg,����`��3y�F�w�Fف&�@XK�"s��f����wh��T�x�>��̌D�/���ΪB <��R
;C�����q��a��~⾛p�>e���~X*8�X�����ZJfN~ʲyJ���C&X�������/bL�ۇ��ؗ8>� ��V���C;1��,�`7��'I��!��&eγ;�`�J;�I���&(��D �k8M��<�(P�;��!6���C����Ì[zZ�+����j?�5c�����^#�L��ȟ:�� Ψ�|J����<2����_ItueY|@�%�I	��ݔ��+���֊��5�&�!�_��2�F�,���'l:���$�K��!�C@$�x[o��Y�Q	�y��|%z��g��
J�6w�R_�$�Q�x����Cm�e�"���NW	Rux�O��.�aTR'SY��֛�0Z�&�q���$o`��'fp�����3�mV��:����p��4��#�	����+rfp�ݳ�zM�NVj;�Q�T<�C:�v_��Jod�,�{J��*�%
����-ʗ��Z�|�!����J=#���J5���h
���L!C���Ld��F�Cib�"B1�C+�c.�b~ٮ��]�������l���!�u�H��{D9m���3|�P���aTΆ��l�|q�P?[��H�z#��ɐ�x���U@�F!Ձf��_�
F���#��kP����Cc_�s𛱯Lc�Fy�{�R��ؗ��V���,ӟ���R���HvK4q��fw��[���t!AV����n��f().W�hP'��N��
O$w��z��t*&��vc��Sv?'���cv^������W�SZ���Dd�	�Q��tD�������^ğ�2�;��>���L�w\����C�*�Dk�>ĩ��d���~�����lC��Ӵ@Xr����"��BQ��y�G�c?�9e��y ���O�@9P��Ǹ�#*:���Y�����+�vH�76V�7�n�z��ԕp�K=�TD�5�f)Κ�"�l��u��O3�Z>+��뺍2����<���Ň��A�������SK����8�Si1��M�Z�#;b `�?l��6�}V��(�6��;o����!r3'Ae��Ҍ�������������Z�eyݼ�����ճ��B�U^�ZA�zz�53u)$�IIˉ�'����+��N��xX,��rU�c����7�p���U��a�E߆z@i���������L�5}���[n����;=Z���J��N~V��\A�!	���FD�I�����`)���G~@Q�
=:�{�Ť���BX<!I��~�~@���%�/�Nc���U���1�4^�hÆ�''�G�U@�.��vX���Ŧ2�m����{������E��f����_ �̻1��h/{Tg$�A�����d�"���+m�/������ue��3@�PZ�� �B@��W��h��Z呲�$�b�.���I04I��=���mWޙ��J��>�}rȊ[9e������2���82�h ""���dH*����e� ���z+?!$���Ţb��*��#?�m�����0�i���3x��+M���c�@��
�,�qD�����{��$�Ս��P,*��?��Ĭ
�'�ϫ�?m)�&W9�QZ׊cy�{��<�+?��!$�|�(��x��D(�T*s��6��=�m���D+y O�X `Ѱ���^eH�A�>DV �}#&)���~}��ɳ�0�fh�S��'��!ʺ�F�נ8�O�Wk�^��x�W>���R�HÓ�A���gp�ϟϒ���z��a���&��,���:i�H��+�6)j�c���3D�����l |݊�$���M��� 1K|q� �Z�f�o�U�@��u�y�T�翷���]��" �q�i�l 3B��-%����<�@Pa��5����&�H�@ �IӜ!�=�Ͳ�#IzBc�ŗ�������!����N ��Ķ�YB@�γ��w�,o\�W>O�SJ�a"��!�`�~7􁬲�'�:H�l֣�sk��8`�i�����Lȇ�}�9gL�cb����s	}σI10��A�J�u�;�IO��D��ph[ϡhz���N��LL L����I���HS���O��nd�x*����&��d��K�*���ش5��+hmY��t���E����Ƶ@M^7���sUI�ٟ�n��8�NJT� va  +n��p�R��qW/���pњA,��k�<Oi�˘+�Đ������`e�º �UM�&�.ӮwrM��a�i������^*�W�q����{wa��Jkq�^��k�f������~W*R=9&��qb)��N1-��[����p,���Yf�ESq���{��}��2�n˓��D�����+Q�R{�z�?����Q�$��́~3V/���y��Q�C�1RT��wNy�߲��s�x��'0F�?X�"��D�����aHD�U-_�y�I��T!_�U�g�D��)����}哅�!&�%�0(l���:�z�1&f�w2r�Q7c[++v�K,��+������C��c��EN̵���p�x�HH����,f���~��RG���p�����o��7�Pop�<vt�?tu�XI�r��h�$�<c�c��b���%��a�'�2GY��g��\�E�:����b+R��r	�s*���6k���J�Q&��Z���'&<�VHP|��ȍ��DHC�&
���1Qo�g� �1�Qa�t�Wr�BRs�o*]�f��1@fL!���)��$��xl�z����FSSU5
�_�j�<�ↈ������7�îJ����7}�.uW�b�Nt��[��7�C�����8��<[�Zd�M^G��#鶙G��nv���EUú#�{l�u�?҆V�Y��I����Q�f��:���R2�)�'� -�`�W
��դ®D�n}$��T��T��5���"�u����L�6C�,��A���5̓/�@�v}������wS�uko�:�}o���G6>,^�U�*�xA+v�(mk�O�lc��� N!#���{��W5�)#����;SF�����ƍ�Ș�(ПPVu�ju��i{��9K���b]�b��̄��S!Ԁ��_:�SK�
�s
�	d�5�K�,Ҟl���
Ȍ����~��U��QրQ��Y�y��0�g� 2�Jƪl��ä�_!�͗6J3��w>���(*Ty<~Mk͈��o-��r���u��J�/�Hl��{�$��� �P4�;Ax��F��QC��7gT@+BpGK��"#{��5���|S��)�!l^"K�N���mV![�$i��>T�+��r�ё�L|�����\w�r�f�Ke�G|Hgg5�{�ءtǢY���_i���W-���O�}[z���{�uϫ ��JKTP=�#��i�������J<���=+�uTs�~�	��9=�͹m��X0���ȿ/�$���LBL<FJ�q\�}��1�L�Z�`HZ�.GK��)�WYy������Y;�~HK�v��x�^�F��(�CqI�ͱS����U>F�N`��9��?�~�07�2ξ`�*P�&=�O�;�cL}ْ�h��,��򢜷�`!	���|$�����m��6f�*9�p(��ŇY��� �(�xs�=�rg#�� ��6�0���)ht*R�<t�dU,��㒎}
�{�	��Wy*�{�f��U]آ�Ւ?�D�nОz�u�0�Y����~D)dAĈ���	�ha&?	I�ê��礀��e���v�a��bƅB�m�Vi��ȣ�T���S$�f$Pf�]�w��䉮����k��nE#@��V�$��i]�Ƣ�N8��K�~�<��z�V��r�J�a������'�#�;�G}��%�pɇe��C�k,��x�Zj��M�*e��X��P��M��Gl���yP�ݯ-��%���z�)Z�; � �&���Mx������+��Kd���#~Y��e���k@6yq+C���&�����&�}�k�"�=�����C���{�R���*5��!~��zߌ�YY����'�7D��.��'�c�5��ڎ�b.����T�j2�d)��-ikb/��8��fX��ݮ+�?1����o���\1��q��|�CN3&��1��%9������
�Y�]:v�BT�:��Nd���$&��=�/������і�� �����7���u͸$!�Q5�]<��Wqa�Ŕp9���(�ԎE���0��:j]M�T�u�� (���}�����?*j)���`�&�;1�6���(Uy���[|qH�T�@Y_�H�gkfn��N����a�z�R�^+����X��S��˕]�YI����|I9O'��j=²c�Ѣ�b@j��f�(�?����0�)�a�$��"��\�$����!�;�i�/.^)eO��u#�L�*�V�������xޔ>U��Ox�(1�>g2�V�8�%rs�6r�gX��P� &w��[��։�Kw��a�!RJ������y�ũ�X]L7�BT닿m�#eE|3tBG���ٍL��oD)�ϑ1e TB�![��I�uU���zq���IQ��y�{���U�����6:/96�[	����y����P�Z;�̨����S瘹9�5�Ԝz�!n-9�A�?2γN\��(����g�l+��2�H9V�����.�!qz��;nA����]��I_.`��)~Р*p���F�hLr���-\(��U �@��[�X� Ű����Pũ�w�ϳ`�d&`P�M�Fyz|u��>;�[��e1��-\��8��CQ��e�1��8�;�s�� �3�=�'lKn(�o�֌(�!'w/�ܮ�Ps�	�H�	lq c��f���������α*��@�v��~��5�<>mT���H	~F�@f(g<4�Ub�8�5��h�'`��I�3�i�E��>V�G�ʴ?�'<��so��'�~�Y�t��W�F��D;�g�9]a���uFn�l��k�S9AL!|���g2�id��>|V#�����k%�Ǳ=�ʀ�GOyb�g�S-�m�bV��yt2b��PR��r���|�!sg�v�{�w�؃�5 �T ��z��Ζ��s�X-B�_ɇҿỲq��R���[jɀu\V(ج$��yT�.B���+��ŉ�^M�[V���o(�y��k[򗣰�:�	��@.�X�@�W`B�_')�'����x;R���Q��`�`'��R��D:��<3Q���P����B.9Ώ�;Z3�ZVx�e�2~����O�;�x� ��Fx��\�/$�e�v�oӈتCtu(���̿�ܗ ㆾoz��J���r���:���Ywۤ`j���;��Z]��z%�y��s��s���H�]�b=|D4��24�d��%SICöV
�(��ƻ�I�s�f��&K��6]C�������ۅC��}��7F�y��!$1�1�|yjoo�4>O隿���ƜH���w��?��*���ԥe{�;r.�@Y��邰蛺��/c�1�SjbO��7��w=�)b��[H7ٱٻx�fj�}�'ҡ&$�ϟctW������n�	�=���8�ӳ,[�9��)x�:�����GCs�J��}���)�hx�%zv��Z^Y�Ry�b<�X����lN�k*vsq�.Q2����/[g���ZF��	@8L���f�V�ը9>R}T���1�d�-�?�����q�K��DI�,�q��3��8�!������_�����t4��iaC�Yd��J�42U��r#y����J��,�2C�U�oXL�%���:9�b{��D�!cqH�̥y�z�g�S7��wxY���_�=�h���3{Vw��CV��U��C�=���+A�܂�`�����[�G�,�.\�b�/Y�j���1�A��OT�bmWf/��;\�đ��>qS��_�k c0�&W�9D��t����[��QQ"g��$T�����I��\#ߕ���8�� ZS�:�"�-�z���$z��O[5���̏��A���t0-2)ȉH����Z�_He�E���Գ��{k� ��
m}@$T��>7$8��T\�P1�%qLێ2��c1�;�+�u�:HsB^��{�K�a�V�Ę���Ô��)��D�
����}i[[j��総=�1����v�@1\��/�������J���QOc��:3���Q��� w	0s���!3���[b�ݧF]�<i��R�=H��ݐj�e0��1 ��r�u}c]��jVz]0����5D�D�:g�k�2��
˝��Cj����`Ϝ�L� �C��,d�:�8�E�!�D�&L���E�=�v���x�l��ŋr�G��v�}f��ېx�1^��:��w�to�I�Bj�'��K���p�����Ϋڸ]�k`��P�/b��Ė5x�����+.`)�^m^ɡ����J��K�9���4��>�W]�"&[X�r����K�׊/��<i�_o�#�|қk�*iɪ<D�)��w���ywŰ�Va��G+�΍�N�~Q����3��7H�fL��9y����F�᧟�1y��S��@v�c��f�<�Mpw��?��\c���a�5�0��]h����	���{0L����5<��sĮb��P~��D�
����2��gV#4�T/�-�wh����Fu}I[-�?�*�����U�����N�h1�_��n�/1��l�`�i��ȊŁ^HZ�;��"g�{�w�/�=��%_.��o2FMP\�Pv^6���&����b���zٹ�1R��H6r����8TdM��ߞ����ˈH�	�>���Ke�#�'�I�G3��r�$mR������7�
L���1�}�{��gG~��O�
�	1X7�x>����I��bH����ҭ�.p��T���غz��Wj���t"fW�с��	�$/\W��ر^����gCܹ��l��Ø�ϙ��އ�l�4�1h5�����|���yU���]���<>�m� �-[���n�1K�*^�䍬_�G�q[O����0	l|~���~	*4�Ng�W��Q �����&x5����Eޔ�Q�`M��h4e��Np`Z&ˀ����Z]�wW.ox��Y7b�=��e�5z�p���(�Z��lA��[��RN��ٜ�P��Hs��I����@�o�'m�)f�
�vcT7���7wԠ��'�!7��x��	�*�<��r-}�zA����jG��x��w����Q�p�y� �#��Q�H�h���>Q���a`O��:�oSC.Q�I�P��*�J�)��V<����;�ٹ��Mf���P5���"�A^��Z6h(�����>���7O�ݤ?�a3�FƏ�W"�0ҵ�)�a���g4<yѸ1�u�75�Ų���i�RW(\�����u�����i����� r[}�1@4��h�,y��I<C�>L@����)9��w�[��[����DD���S��J�(�����'���BZ/��c� q��x��4���X~('��X�?MF�O�z�[#�k�Tv�5������b�㴂8F�|���P��s�?��SAD�N�@��F+��m��?-������)hi���X�������Ê��ş����j�b��{)4Ddy�ae��p�1�υ��� �%�=�0BuX���!��4H��F&�bq���Pĕ�g/ITs��E����尾��Ч��X�dD�gL�� ���[��VZ8]w�σ޲H�s�(�Y�!	�����%�4��+�F~S/׉ۇ-�
u�|j�"̂�� *$�t��E� �d��3*�R:S�X2���������z�s%�?��*f-6�U�G�)Nx8b��RPZRbxܧ��3R}9�w=c�'s�[V�J3z8��!6�sK����D���ƲFs�CJB�Qٗlf<K#@F[��ZDl�Z�T:{���5:��I��=�G$ވ�����kR0/##��%��� d#-e(3���.������I[S�P�Xr�9u��h��
�kZ����Jt�ץR�d��My�Yˬj��d��&t�1��s�1�x�B3���zC�p{��]Z�EX��z�i�Z�J=~jM����%)#�3�qe�$��j��0vOM'�+�;GҪ��@tbL��~ʶ��V�^Iqr�˵!��u����0߶bX�5t'J#��^��}~�/��[�Ős��Ċ��%�����_���@ᤆ��^�U������6m��%�f�A�0�
@��3Y���e7/�gn�\�޲��:�5C��|R���I��zyn��J�]�B�'p�c��J�%k?<t��d�5�i�2��~�����1�gY|G@.��D�V!H���h���������a]��!C"Pm�Bܧ�5'r�k�oR=
eƤ�z��E�Nm��^h�R6�Y�wr{B�c�zÙ�����k�M�T?6>�(X��#֝K��d3;�90p��X
���P��w¨~�טH�J*s� Ϫ�W7�qV����j,��d�e��,E�7ƙ��Ƴ��0��U�[�2�@�VQ� �W`�P��fȦ|��fKGED�5�ao��-�_5e�����34���Ǎ�/��Lb���Ds� �:]U ,���2�?��i��w�� Л�z�@l��򤵛ǔ��z�ǩ4���?��GhI�!�L�Ls�g�h�pU|LS���7���iP��K��|���c	��2v�4t�f�����k������A�fX����	WH��Xɿ!�U��]p\�M�W���g�s0��u��%�O���6f�4�ZPPZ#~�3�H���� �������#+��Ճ.k��^�V/���Y?�K6��������<TA2�jɩ���VUQ��b�Ǹ�w�/��"��y+��We�m}��3�M0�D�V�#�����|�+K�>mk���tmqO���0ơF=�y�i<��Օ��K�F	���37ۻ~�D�A{����,�'�� (��d׾�ZNg�������C��I�QC^�V�/yZ�����6e�+!e��h�U�0Ѐb+p��	`="�l]j�Kb#W�� ��ܲ�f��j���e��j�>?�+���Yrm��Y$l�ޖ#=Z��c
r>Eq��K�q���V����R#��ec~dA'g�V�,��d8���j;k��� %���Z����=d��|h@�\���o��00"N��?��cߔ��x�O:�� �p(p�QN��K�G��,B��,[�m
4S��ak�D��B��;��3$�};3�+��uJ,?h@�(4������>���)���} ��v���%�3�성}T����K�:����X��|����p�v���fʆcOD��ҙ�!^�OY\ac ���b���ݸȿ3e=�hh�I�h�yeX^˔<��$ؤM���L�7�^���^}Dּ�,�r�@⼂�.	2�*!$�o���9�����	��slw>�+�hP#��Gp���,�Cuކ��%����R�,wo]h���.�W��P�Ҭ~�n1
W%	�| (j���P�����I)h�J���������7��c�rF���-��оQ�P�s�����/��l��&�a�H]��P��[BϏC�_��~��c�s|]�/s_�ɢ���r��s�v�&�F|���*1 n�a�j�����$O֓���	\Õ�6��f�bՃE@����@}ndpr�G3ȴH���')ǧ�\H1�a�����u�:��>�Ƹ�LuO�)���-
���t;���$�E��l�=��8A<��|�t9uj���>B���>���;�'�a�b��Q!|�t�E�e!��2]�O�*n���T���6��t�ǝs8���!k���� ���^�)���|��½�\LI�c��A��c`�f�u=�� �0Y{^$��Gg�gY��>-�L?�w�G�Q�[y~	����L2�*�l���)��ta��kt����[�RA��H/<w0��~��e�rt�i�t�x��66��دl���?č��[^0����	�S��P��q���N������|���8T�w H?�ʭ2K�[�k�q�5վr��g�e�0��Tc0]�>	�kKC�n�c;��
�t :s�~3En���c��6,�9���x�M�KY�e�6�c돲{��H�H�STt�o���	��qe�(���T��g%H��c��*Յl��·���chr�x�²�zՀOr�e׈ll�nPZ�X׻���A��ɼ��(�rx�Lx�9���@!_2�E-z⋜��u��e�/׸�Rj ���~�:�ݤ:FN�i?�nH4�t0�N���z�� �Q�p?�z{����-���.V�/6�N�^>����w�-#�E}�����p���n�*;S��IM'�t����tS�D��kr�!�=
vICd����%��Va�u~�Y0z'���c4�U-3�"��]VhNS��f����s�94��DN���W���F�@z*�V���p>�u��I;�^�Z(MY@��PξM�0;� _�W�Q�j�~�+���0��X������.%�7����t�W7ߢ�?䃷��hM��(�V� �7N��O��x�}�!)^�Q��8ya���6�j=���3Q���`�2�C/@����ia��P������p�~�FZ�l H7ۥY���m�|��;���\g�v�v�|��}��Ɨ�g�ɧ��8�����G0��ޜ	^��	��^<�(m$%��8�ˑ�o̓k��`�����L��tc����R_@O'�7x1�U���U���C���$  P�)��uS��5�ț�W &�uukq�W<`�z{��%�{.s��C�3����������q���[N����7.=7ke< d]�k�8�	��Q[�(���f*��AI�C�(�^5̚(M��k�cԫamw��i�g��t�k��<��ܪV��d�]�kK�8-j���K  ��[:Z�8�1�&��H9X����4#���Q��q�r��3O�Ndn��ጟ�\�Bǣ�z�T袨хq�,���F�ov��H�Ck���oU��'��1���.D��)һ����ǦnŅ��Wp
>�
�'b�}F_�o�����ETC�ٯ�$*���&��lƬ�j�y��\�-F�(!NeF����N��|�n�Q>p-|Of6|g�;&Y�H��i[�mݭ��m!_�������8=:��*d�1f��Ñ�	���>�W�yۡ1��d�Խ|!��e���ucAO=���=��Uv�rTo�`ȟ}i�+?��1�x���b�	3��v�.�Δ2��~�x
c�>'n���p��P��,�q�w��"vr�Ìw^ �9�*օ�U�~^�+	R-\��h4�� �E唉�$tC�3���(����ؒR֓~� ��=�H����}m!��Vx�xi},i�wO��RK����fV)��1$�R�P멜w^b7M8GJ�X5rs<a
�S@.�Ia�f�p��#� N�^R� �T"Z�A/ٞ�p#/�!4��z�L�(x.��f���&$D���&'��A���.0lK�f�ISލ����e̥�3TV$t����S���ߌ��gI�Lo��w��"7������*��Y3��jHr�DBqEcg!`Ks�ePIil���y�(^�}�^�T�_����d0�����n�$k
�� D�u��˘W�ѿ���2��5�A��y(�Ŕ��	(ܾ���k�{xI���>���-�=b��p;�|9{���z��J��``���5*m*��"E1��&�ʠ�{c�`v�3h���F���q0���z8�W-�7i�=z	շr��C_L�ި/q��৆�l���K��:unz�T�W���x��+db����}��K]����S>�|�����3�@p����˞�/n�J��]Ů�Ȃ�\��ِjy�P=�u�Ɛ�+����m�i���L�b#������G�i���M"�}�8�Ĥ�|�󁳶�Y�0|�z�f���Xxѽ��,�˘*?������q܅�f@�L$r��Yt�A�]�ŶC:R�#� �쁺s�1��Ԇ0��t*H�0�B1��*�4�	�P��F�Ao:v\�kCB>���-�ԩ��:"���>�C>�ACdvF�;�Fkv���QJ6;7����UI�iO�3(���q�K��M�!�v�(��դ܋��Y[���aw�h;4�LvoQv���`�.4�$LP���L 28n/�Ƹ*eL�zt��f�5�R淮�ӥ�+��
sϜpdڟO+�S/2��Wƥlm������WL%V����=�/O�!ߠ��Czv8CX&m����/�/���k�+[�Z�1�Kn��g�|?����z�F�Z�͸�YU�4���_��dx� �d2� :m3�у
�e i��)^���O��.3�x�U�4oY�I'��0�(�c����a>�t��u�ȴ_9E�,>�S����:��!��{ҐX�G�kXTZ�G:��k4���|f�B�����7q�u��jfR�L�ϡ�Қ��C2��D���D$L�o���:�ՅRomq�.	�T�RϜp�yZ��rP��j�!������P��}���.J��3�.d�>F넞�qZ�s���������YV���OD���;��4����y���|��֖03��r}H�!"nߺbG��	����?�#�Ȗ�H ��@�χ"2[W���s�4�
�P���i6�?�;�����h�O�#�|>%��k��Jh��0�3���2�~�+�d�W��3��.ө2����p�@��c���O/��6�dk���-�]�7���y@ks��חPVwFLRL`Ic�^M� ��xjX;1ӎuh�U���yo�|{b	Ju~8���.�����RX�H���"��^Iג�񄲚��J�t47�(\�}l�d>��Q�y4 {�aڐ�i�S�����p�'�j��@t^z�o��df�Ϥ$V*޼����9癤Tg�������	䐷�[�"�r�PM�p7�8UP��>�d����<ݟ4��H�Ɩ��+E[|Ƕ�����
2b�����\+}��MN0�)8�w���C?6�L
�2�gD�Y+?@`-����Vu/�v�.ݩ �oL�9Q��׼����UeP^�P�N ><Ѳ��wÜG<����O�D�����<o��iU���@X}[w�#�^�4����� ��s�ک�SY����ϧn��3�=ѹ�
6�>�����FZD���R_i�-O�+k�$4(_iu}h47�0q(śNߡ
G�A�a�qX��=N�� �`�F/�!x=\S�7#~g��`�g�1���i�ڧ���9(��p��Af�FF��/�kr,\Sb����a?*�¹��x�O������ҟO�;ɾ��p��1��ҿ7��Ej�	�>P���v\��I�f�^�A�I�����ء��{�fKm��u����׫�� ���V��B���K�f&���>�Pk��h���Q���@Z4��)����ˇ�ko�Mެ���7����W�ެ/��7��~��u�5���b5Q0y�Ig��Ib�jB�T8��g^�t�D���^��Kv$�O^��Ns<KWkx<	�<Dj̱ ��,p��P�"�*ۯ!�w���'���}EOX�np��N�Q�.W���W���!�_��l\jg�����X�
s�.|����}Qʻ�gJ=r�T���S��jG��~6��&�&,˞*�>r�:�ive��KR9�v�w�.s�y�NbX�kN�rP������@-4@�3\�b~�3[�QF����a���M�i�mv*@M����m�_D�6�}W}���I�=�������e0�L�N�_D��5f�%�v��O����Ԅ,ڈ�n��/ky���(���c��y=J{<��ѕ���#ag���8�M�����ĭ�a�'�o���a�ń&��;-�TQ�2�Ͻ�Pj�Q>����mmb��R���O��$h��_�Q}� $d�o8zm�q���f���n @j-dbl��ouM8A46'����<�k����Y�k�-)o���]��6��]��E���̈�	ʑ 0���]"���u��$�����W���>�`eG�����>5��"w������!a-��E˄�!�� $Xe�Y$�E��F
�Z������0J�v6��Z �& E����[�M���{�6W��	_�ʶ�	U%D�5�	J��.�׭�Ds��U�����d��q���1h�W����5������aD��e6�r��g�z ӹ��@�	�0峚Ϻx�|���\��3i�Z�0lK'P��3Q��t����k�a\��9�7�k��z�LǞ����o*��J�����~��y���9j6�_�Ι���/�t�8�ͩ���8Ú��0靭{�ɫHz��bsg�EH�O�e t��m�0�2+�u@w��N#�4���Om��
�G=�H��y�kN�8�P"@#w3o���U� XƢ���9{]F��h,���{���fg�׆W7�s����چ'RW�l�r��.m�G���ws�ow���Q����U�i����!V�5�iu^��L�<�hG|a~���)ʨ��������F�1���:9���FL�w��w��^��)�>bA���<�p�rսspfzQ �)P S5��#Xm�&�3"�2�@���5�r,+Sｶ�
��v��mS_hf�pu�Vv�E(��^/�u������Р$���:�*�A���F��q(���?�?C���<!��	9��Rvz�mŸ~΍9���OH�"�������g6,t�8]�gF�*�*��~���>-������#$���N;�ӯB�Dj?񡼇��/cC�a3��R���m$��0��Эa�ݍ�����Z\	��{l�@Hug�kU'M�����>Q�3[Zb�_x��uSy��8?��#��gH�r�b�-����.����C��"(���b,yǢ6�#�[�Iφ�1ߑu�R5æժ%�7"f4�q[�EI�#���T���t׻�]����O������-�z�E8���K�j]fF���5Ymu�\�ih�p��,K�SL���l�o�1���}�x���(&��Q�߱�e��׸A��*����#yC<�D#�]w�\r�;�Am��3��>]^kI1L�4� ���<7֞7���*ؤ��`�~|!0��^��8P���# +��*�6iꖆ6�W��=H�ba��`���P���ksh�ĝ����<䙒:�*-�o�VX�Z��=�B�J˭t].oe���O�٢"�����ӡ2i®SId�G�s����R����A�h��L]���HE�����ys ���+� �pt�F���R����3����)ˌ�X1N������q������g�p��3J�M�� {�����{e�rp?Z`E �ZهtC��R��&b���p�vG��r��#�//�i���tI�z)���]n���@�Q�%�<g���<�H�M��o_[ܲ �i{&��7�Jx��+,�^5���ӸP�ۍ�;k��9���2�5����G,���2��(TJ-OL�?OnX^��I��b&�_G{`��Iʚ-9�0��bf:������gڴ���_4 4+����:�2=i��qN��i�vjy���L���ݺ��"��k�ԁ�U�^,zT�7l��&�B�e�RZ~����ay8i��Bʔl�\�(��^�.��$(>�~�!��ۇ���H!ҁ����H�ᥧ�����K�}yXїjU�E��㓅_����e��py����(��z|�j�+x�����m)�������Oeǖ����oY尽��k�n���d�� %cE���y>����4e��@���������t"����$�"P�u�+$�pS�YpQi[�X��r& �Ի��!���m�4�|�`���15$Y�8|FJ��j0no-1Bo�r��}	��a��NA��p!MT  ���S�:��+ѷ�<m�(��T������j����������<�k�e� �ސ�v��I2Gֺ���Dw�N�ۢ�$E����p�~���'`��� o����o�/l��$-�F�b�/~Ur^�f��X�6��8��� <&m	�Ec����y�9#���N"ג�u)4�sBʗ�F��N�XF�I��M���o`ZC>�B��R#��)
�� _�	
��=٣|B�3w�e���k��+���JVQ����v�5Y(����Z�䄍��Z\L<tM-{��E��V	��f���Bv�O�T�b�|�G�~"d��fy����F�[<�Y�Æ��q�ϒY�g�II������b����05����ѫTh� ^E��&����]4oeǠV��&u;�_��q���E�A;z�n"0��q������0\�M�h�+���4��bC7��Ю�A��.����C=��h�b�u���p��{�V]�L�%��(�_7gk�&_�d��t��N���ť��d>���kc�["��C�и!�w�Z9~���]�@I�k���lf%�X��j��� �A�(I&;�������D6!��Y���O��8�o+A5��O������6��k�^����(�� ;
�AZ�"��1f
Q�4���Dk92~b�,bYH?~ZU(Dh4}�pZ ���������|�v��3���Δ��bt���}��lҌ�;��7bi ���q������Ռ�$��ɛ��S��U�@�~Gm4�_|�Ĕ��������p�P�Z�� U��n��gnw:cD$ �9B��h��t����~{њw�B�5&W��7w<��%g��6u7�~a06o>0�ޗ�PhKT�`�2Z+?[ �������2��0O�*���J�U�/q>꧇XI^��,�K(;F�]-���5��Pl2�DF ��� eP�A�qƟ�3G�����P*	(�Li�:dl����=���p�=���^�p��v��c&ur��^̦Ƽ1���>�
rH�N0��M�A�C�����F3斻S���;�D�n��.V 3̯�S8;�?�-Y�M�&�E?�����b�.)41K�I�g@ac��dk`'(,!�����|��ǯX��� ف�]�}��1u~5^�`�&T܇��Kw�rkUҘr��1P$�9C`nG܇����h��j�|� ���_�Dgd)��:�1$��=�U���)�����_Y��xЀxi��$a0=!mLq˲�%�L�?ǟi!�A������wD4�<���~�k��xE-��Iy/���أ��Li�ו����h�@��0]E���tBhQ^|7��M�T?���@�ߵ��/���U�@ɑH���cBdb�Б��#���k�h"�Tu�1De*�s�7i͘0�_�~V
�T���R����M�¨���l� �^�]�W�-��u���8��$���#c�jj�c���\V�t��O��e���ѡ+�����*+�4PI����)n��$��Mv�\���U �k83	H��1�"
����5��yO�D�Y�=���R��F�â�غf.��SF�������1�~ɍ��NH�RT�]F�:^��ay�~�����@��
�f��Zt.��!��ܽI����sz����9v�7���)�I��k�u$�|��݄%\,β:��(T���m�mC��z�ÖC��6zI�B��z��*���N���m���	C��y���>�c�L߰�1'�Y�_ۦIo��[j��܏�xC(I2�����e�̜> k�qM�ʕ���c�0�v������y��<i�)��7H��t��bW���zձ��w�������Mf�X���p�,��!�T"�7i�����E
�^#[��<�9� ����%
w�-C������"���NQC�͛`�{��}��٥Ժ��W{xT����hCd�0|��n!�?�f�}��/v|����&7lZu�T,$G�ښB*���]=̀�}�ڵu��v��E�Z�[YS�w%`kV��4C���;Qig�;���2J!{?�L�0�'�y�2 ob��G�v��HM��2h�56m�ti��AR�֙��|p�x�d��-_;\o��q�����|��m�:N@P�`�������g�QF���_=vn�\�7�hȯ�Nv�<B�A��/���,0�[	��� ��D�X�i�x�M���2�_�F��"D�1��E>xv6���?�$g���waf��sa���V�0�����$ϰ�j:�U�|������*ês�X��+��
���mZ�;����MC��>̺����9mw��m�'�"�En��n
j�(Е"ySA@�9-�Nn	WlJ���߾ ���,1]�a��@<�x��<�g��͍|���}�9-w��� E�f�
��P!s|I�w6�_i��؊;�foK#)�����x�&�)'薴k�YU���˥���֣�)ꎡ�B�qd�,�����[���9��iW�϶�d�C6�L��D^�&k���7�9xZ�X��K*��dA��*�v&�M�K����h���	����!�Y�8�T:Em��6�0�$5��V��W�����$+b�v	м9�Р�d����ڷ�s�����vg�Na�C�����C0��i�DR\��A@"�?�I��H�7e�ԑg
6�O�k��#��u�����A�?F�2�YX�y��
R	N��*�?'_?�R�^�,b��O�ɽunJ�#�7���~D*�A��=��:.����(��lg��zԦE�Z�j���EK��=E�pD	�0;�o���5,�H�;�E�pL>�Ү��P؁�T�l �O�y2H���u]��I$`'��8^ccW�>�L��.ʅ�f�a���7#�&����_a�/�/��aSZ���zlܥ��MX~��jO5���S'�#X�~�vѨ ���z�G��	/��"��QVP�7yq��{�
k�0X���|s�������iCk�X�R�����q�H�[<�u
`�F������$�窔�W�y�@���]�<b%QN@���k�����t6��gMH�T0����I:�9N��P�B�O>�u)�t@�đ�.�!8ŵ�ᘨ���\1���"��(�c�^�m�?"L��:D�:P����e��L}�Ex�$��� D��M��Qq �g��2X��o��J��}/���|\R��������I���ۑ�fW|�oXL�U��Ceĉ��x�!�e=�����
�b��X���YN$t�{OA�ܞ�O��t��G�/���5���������o. �5��Ň�B�ol�)������0{,7�gP�>���E�����MU�7��Ou�J�J��]Hd�Ϳ��O���.��H��H�C+�ML1H�+z���/�My�$YqLg�eWg��2�o��9M��3��<+X�����T�,�Q�5͹XV
D�/�lp��v�둛�ig`}(��@���B����k����wG�e��r��B(��8�x���� ��WB���1_|�_�Q�q�C�(KK��ds`L�bBe
����{t$j>�� vW���4|�r���h� �YI[��Ɉ�_��PmPD��/�L�=���pJ�j�J�(Z_����q;��p�@�A�A���r��6\?Y,*� ����2&φ|@>)���&�9axd�^E�鳄�t������81�+@窒�]=�E$7^?���5�o��K�B�r�A��m�4u01���y�e��g;"�MFĔ���èv>g���򖍬}�`+�ȅ���ji�}b�g0�*F�C�����"���`�ݖ�ґ�^2�,]gͼ�4�	�/�w/�ڶ���|�F?h~����ו\Y�eGf;ٜ�ʟu�Jw>`�G/�r	�t*dq�-��Ɠ5����\p�y���Ӡ��D!t0	�7���>��L$��?��P�E�'bb8�瀝�$�8��WyH�K�l��h<#L@X'���?��-�[��W��2�+�[�̫�$[�s�6�)׬�s~�{1B�D�,���/F;%
���g�D��Cy�Ƹ[�v+-.ųf��}����@Y�e�p�����[]�3��*�֓W0�t���*0�k4��2bd�;�xᆛ�'�g�c����N��A�(Z��=�H��VK�k���'0:�X⬆g�|�k'�/w!���B4EQ��
�&�M�LkU��s�X��֬t�.�wH���v��.A�s{/���I�EdT	�Cj���Ni�+EO)\w��2 �ƞ�4E��
g�p���L�H�����Q�|Ɂ�B宿�X�{#����#��
Lm�u84�,�e�/^�ݱn���@\�����~B�>�T�no.D��(6����؍5v$M��6T�x.;�rf�я.�i���s}�!�����_�V|q�:Ϋ��?鹘V����ϙ�1�S΁-�}Z���(Qc��F^��3�<�w\ue�R?tb I�Z1�<N�E�v�0�i ^��P3'#��bXMN|5���������e�2̕��_p_'�C��4�j�`�W��6���J�uf�>���jy��恓�e�ݩ$��4-H("�*Ġ�Dl'/����ED�:�n<��<rn(h��~6��H^	C�&:�:%���L�S`YW�wB���e0�ZyÞ��R��X0H��KV-٦<F�~P6�po���.�r�����7�=B��|�L�JW��]����O�����8�B��3۫�z��L~z1��"�;ȼreB�e���r�����%!��
�Q'�A�@}�����
�c|'���Y�#��|N{4�ϑ~XI8F�`T�v�fu�n��l�-&����9f��5��c� q�	΄)1Hn�o�ǲ2�>�M��Sh/7�"��B	|�}2�Hǲ��S/�
�h:�C���A~�?�]��Hjϭ��K�)O�7^�$'����z��3�j��^�q[���8�a��a�����Xo
�+���|R!�EK�׶ޔ�'Tt�KSM��q�����B-��NA/aUjQ��i"mP���h� �� Ϛi4�x~"6*���8un�<���깥̈�TOTL��P����.$���"f�6�-Jp��Z�,�~8#=���k8ȯšPא{�������R�O�t�>9S(	�
�8j�Ꝁ���:��r|i��٤'#gؑ%��\�)�"����x���9�(Y����U	8^l��U������/�6d+�)�.Er������m*� �Y7�X��]}ԨZ������%Rr��h�
p��U^9�/L;T����s;yZ�a�3����n���R�qg�q�4g�֕��f\��v������lb=�<b�����U�TIf��o�hb�#hLd����
>Α���ru3M޺K�Ep)���:�~*>�J�솱�J?.y���@S�$�#���X*Mi�ђ�<[}�E2��K�z��t�_Ad9������;!���ܶ�&�5S�<�k���XY�u�����}4���GK��T :.tG�gQ�mrivLC�ewZp�����*��v��$��T�_LcG��ݐ���D���r,��*/\i�����N(�d@�wO ��Z� ��hj��n��/�?��=�x"9pH���l�T�W��/>[����gq������^�|Rb߽��H���2�]�ݣn���|��G}�J�N1J�z�>�L�觼�FZյ���)yo"�,)1��(b"��H)ϡ�nV�ݷWr���at�~�7	��MBw�`�2�п>��h���lQ� $h��1�p{���{Efc��L;,u�C��ܺ�l���^w���+)�/�����D3z�7%&��t1��	bq�Ju���04լ��M�d���z����|h�Ѱ+'07��jjJ3����-�����������D��Qi\Z����,��M��^�g�a"].rYP7W��:C�\r��8��*AmQ�-7�I�5uf�'�����,\� �m,��A�k.�(�O��%\��~�u�N�J9"�;HU7�.n.n��I�l�^���s����V�X���
踓�(�zm�)7� �	��)�Hm1sth�s�`�������D@��<K���8��co�&e%�_Y��Αʏ��E��h�	���/�T_D"�lH�J2!�Ꮺ#Ԭ]����> v�U�a���9VTS7�O44v�K����,~G�	Ql�8t�U,%�����5���5ay���Y�p��5X<���9��X�j����)���o����g�s�g���&)pC2wQ����;���z��CF�Gr�Q�O���t�Ͷ��"����'�N��PfYLZxc59_hj���'|����Ͳw]�?��5ҹ��M��ŭ��zg���S7����OJ�ݷ�;]�Sʏm��1O���V#02�&���/n�!s��!h7�(e����9V"�Χל�+	[����'渢�4�>��Q���v<�$-��:w\&���W=�d���3���h��X��(�($�N~1���UQLΖ1��O��p�6�t�0BJ�K�(���~��~J[mQ��M|����2-k^/O��o��\4ʫq����qv���`R/u&ſ3�+�����2b\ ���&�:\��B�mv4��~T�x��n9�@������$<4\�*+�����nV���5"���)M�gۻN7�G�;`��Nkn���Ғ#���-���{���v쏲f�DYm7r2�S`"��FR�_lNg����:X�8�H������݅a��M�e��{]��s��1]�-4	u�-�F��d7Jr՜:��c R�M�.�@М���艟�I�֩����=�i0����f_��m`�Z��"M�ј�m�TZÕ�
$C��>%��{��]�O��8�fK ��c�R�IkI���t����>��?<Cಈl$�kU&qk��v����X��}༔g��[�k3�����*�-0��&�D�R�m��}��9�Y_��s��zê(ƺV�x8�-��[�_wt� Y���r�^n������ZN��x=9�_z�:+\�_�p��E��9��y��o�m��UR'�y�Gu�q_dƹ,8W�_d,HaV]��m���ɹ�MW�]�h<�kǏ���yB��~I2�\���!��'�&m�v�[Y��~��vD�; -�5\����*�uò����\>(g�;�uN��=����X%O����p<Tr�oa�0/	ށn���,|�L=[��) ¶^~5Js��l[!$I��ESԟ@̓/}��Y��Q�QY��o
A]��;�����W]�@+2:�|e9����@�R��*�B��^C.���U%n��d�"�:SSZzP��A�2CW�p�
OmS�����6ŧssV	�̻��\�lVali-Ď����h㿨�=�5@���s� �B�.j�zn�t2�p������g�Bq��ߑ����sr��m��'&V��?� ���
��W�v,K�G≖���^zK�LV
aؽ�s��I��A}�Z���0����5?��G~�UG�~m�@�$+	 `Sy�J��]=��6���p�Oʨ�"a��x;����\s���N���AF&�Ku���׷"R��T���r]�>�aڱ�$q�G�/!��@(��Ԣ`Oəe�n�s���6a����6��W���e*��}rQ=�������Ӟ�2�_{�@"p��3�����+"&55������&V��<��H'��|G�1��f�`�W-fe�EB[�'(��}�Um������IK���j���iU�Ƽ/��vI���m
O+�K��:���[9~2ç��_[��GY�В�Ɵ��ęB������e�06i����Y4=p��ɹ�SkI��W�����b�{���l�Y-��
���䘦�=o3_������	�KR�*,����2�����M��t����N]E~Z�a��;b�p��#���זYn�>_E��3�ۣ���."7%�S���3V�BP�K��`���{l��r5���ʃ`��xp������uGT��E�t�y��ݞ/7b�97d=� (SK6�K��$HS&���,�|Q�e�Ά���R�D�01d��T���Z�U��$%�>o���doFQU��v��zoT�9~�KC_�`�mh�(Q'y�АV��F�H��Л��^J<����H!oރbE�'`s�y��e�ϗP�aF۹v1�����b~�u>����6)E���%/��g$�i�
&��_f��X��G��,�W��9��'�����T~m�����[W�[������eBϰȞ�c�_�N��l>@�Q���0j�N�t1S�o֛���+�_sIޕ�L��&-�Hɢ(B>�AϾ�,�f�Lp���b��{��\��9P�N�`�<��s&r��)(o8�S�Q����y���?�%��C�H��y�����7c?�S?����G�>���ɔ��hxԕ��ʞ-�eJbMx.V��ȝ�v�bR����0@\;���84��2Ԉ?�+6>��mwk�c�x�q�{a�v/^"�J�J���2nZU�u)̗�5�p�!_u�X��!�F�A�l�		�TW���DR~�J�;��2|߃A2�rR<�Vn�Q.K��́���x�t�؏Gb�w�
z�#F������7-�V._��R)�g���fQSP��yT�W��8�A��|X�������/0&tz�E�hbd��N��~U��r�Rd�{��Q�4�X�#gϻ�H��+$X��f�s�/���Vn���5�ulnE����	�������%��xYH��h)) ݯ%F`��v�]�Y=�������uV�C�1��� �cm�z`��/��$��u�"��/	*��]��-Y����VĒ��FW��ͬ�|2
	8p���Q�S%]�|H����?�ä��J���k�������a�/c�+J��0��������P�b�����gDD�!���M}��3>`�4�5f���1��d���=� L�����������VFЃ,���t�ww=��P�9���O|����|����fwJ�Oķ'����H�س�ea�i��w)1�[휥 �7G�ь��3�m�K^G\����"�Ou��
�ٓ/<(�,V�^ԙS5Bu�j�����%���k�!��;2��]�`�f!/���%�t��a�'�J�ı���L��I�o��U�^�F��� ���w�(Z~�>��#��?82��AHI�p���e�=����G�#H�Z1;|AO]�n�`�®f��e͓FE�ϒ��~����A�}�Z&m���$��yL����t��"��H4Lۙ�
aޅ��dzղ�Y�^��bՂV
���A5�2���������xC�άm��8��j]3e^AǑ����Q��	l�ݛ��)��>`b��i�'?hhKo�Z�"���3E��s��Obgy%�+?:�h���j����1������P ���[��Q��fE���/p�1�
5_��h����Ȕ��
:�S*zԮk�Ӈ�f3,{;p�%�NU�`�P��uc�>de��7( �����d�d��
n5h��-�׉⅋���i�-|S�f\Q�U��lAXo@��/�""?6�.nXωG�Wl�3څ�����B�f��Z�)@���v4:u�%(��;�9A�wy���#4v�zF��{�j�x�^e��ʴԯum�G4R�����U�xL=�۟kׁ�j2g4==w�9%���� �#�k� �j���	z��u��75!]9�Ea�MWX�4k�*��2uF�~Ɇ#�	㥬}+���}�N_��/��x\���x�H�i���EQ�"5���}�,Ngz�S�ΰ�]��e^;�3z�1�Ͷ
��
���w�|KR�J�k	h�{���y��7�ŷ�-\��_!&~V�2��M��&������Aqd��|�$�5������#L�P�������EY��ޒ�Y��
���<FST�YǺ�1�����fZ��>;d]�_�t�4{���g�()�Jw@Нq���#�d�fn�/od5�D�m��V��sȒ Mn)���Kffh�f���}�q�8�6�P1�H���\ �  �МK��B�;�C+o	8�r��,4&�!���o?7�:a;���c�@2eV���!�<�����ԋdbv�{��:��&Ȼ��rKT(�t�R!��(��y޸�b^����P^�0�/��ݷ�DX�O��/Hv�P>�)f�Ŋ�uSެ8W �T��,�Oɥ0��g�>2e���˂"��ۄ��>L�x@t���? ї�d���i�Z[Y��r^I��ǲ���q��`2W�p�~M�ڔ�>f���:�>9��&P%�#���S�u2�R���=�u�@���o�T��ѿy�w���	*�6���E&r4+.l$���
��߈<dW�y�y����a���Q�@�h�g%�l&���q�	��������,%�t�!��#��N�F���W�B�nh��HQ$\��!�P�����=C��~$,Д�i-O��0�칷���0�Pѿj\��~x]�I�zN3Jg e�i=���]|t�G��g���V�ȕdg3^�Ȑ=;l!���ǁ��Q{P�i}4�< s���U���^	y�E�_��!�h��ce[�J�sy�|��fKq�u�ī��;ARm�6�c�q�c(ַ*��`[�{��*�n�ܛ�c�M���C�@�j[�+>��AGMS�
���)��JS�&7?����sr�[[�����4�W��� �/%��oF��+DU���rO�D.�-W-�W�RnΗ���}�;�����29�.�q'ω���!���rѸ�.lY� �PΕe�D���}��h���2���^���	��W���1P/?��E�2!�P�g����St�(�NH\�8j���}�r[��h�Ϩ����F��1(�CM�t�'?ЕW#����|��jV�w 6�`�Z>�~O�~N����`R\����$^���?BH�?�s�j𲎢c�sy��v��������L���P���K�=�U��Eя�_��
:;�$aA/d|j�f�ͫ4t��x�qfS���C%�:���jf�{�!Z��%He��(�0�k�n�ƃ�pU|�q����#�̈�� '�gi�+��ΕDw���ۯ��w�^��#�E&��G	�ff
�'ld���βD�"��O��0��ϖ@���щ rrQ��m3N��;ҥ��B�T��wb�\�YЏ鱆>h��A�����mI��ϧb%�G�l���j����iS ���i��
�F*g�]4(
������:�4*����o�d��ӅN�VC�eҌuJ$\	 �Z��"b��ĬT\�IP�̓��A�t1�dr1�ܣ8����w���ǰ��R:���Bل��_i�*%�Ω�E�9�D�83eoyIU��K�Td���F��i�dU���Z��(<(��լ���8j�� ��Zn<�lBX�ų�N�Y��T�3�"'�&�q�1OJ��[�����^f%@n�T,k5vqm��^;	��j%8�OB�?��-�����Y4� �{����T���tq�8W�,
�J'��D�`�i+����.,�H:���X�'� ECG���G�^�`��j�uKw�1�����~98�n�}>r�����c�8�l�|xQ�b�0�f	T��~�v��Y�K_�KE��_��l�q��l�H=�&5تP�o�ޡi�b�,�S��G^�jj�y��(�������3��~��?��}j,�,��J�P�B��
�q�U��1��tzJc����|���~?�v&�
���se=��a˾~��d�<����e��ܠU�df��X�����L`��'�G�֕v�\6r0�@�	>>���³S2�o�"б[.~��B&��K�� ����FN�5�u��/�e�,��E��C����`*�=�<2��E&@@�����v�S��XI��� �y��`���7Kg���m.�\o��	J��Ϊ�]�
*y `����Ő��%�;�`�c|rj$�W��^���cUnTE�\�:�r �2��H��^���]1�%��;�QAXh~��ɼ̑�EgC ���l��q�<��[OJFӍl�E�����Y�8ش�E��'��w��O���>��h��<�������Mֳ��6�OC�9��E8§Uc��!g��0"��CXVK=oġ�$;%�c��m����� 'U�ڵ����>��(ػ15-��oͨ}��c·���L����q��_�@��0�G�q�ޒʰWX�Ba�� [�דr�7gNϰ�{H���r��Y� !�`;�����ɒ6�;�P-w�:ai8=��6�V�	su�vp�u[��g����g�H;B�� oW����>�C�e-?����0&}
����Ƿ�4s.�L蚅������?8�{Ӯ+ڊ$n�88[����#O���<!��V�)�t��J� w��м�Z',���a����^�-ۑE67�M��C�^=��M)��D�%t�ViC!��nhU�xZ�!��k���a��׫���*�����ظ����/Ա|@ ˭����RUճ��G����y��:�Aԉ����+�{(��H��B���4��eX�F e�c(�l�^���8�,�t���e�U~t2��^�$$"[��,r#���=�:���Q�HLw>�%Z�͵����$���&<�#nJ[��?Z�~���P�g3�c�C�
�����U?��Y��ʹ�r�2fx N��N+N�Qűo��q�����_�"J��ׯ�\W��zH����Xݶ��8�Z�_n��&\��Kze��Ĕ��X/�R:��Z�����0��X<Û���`�j��3��>u$bM�`�3�Kv�H�p�Ztm���aC�nW�,���'%.	�k�c/�Z�(@zy�⽛ᶤ���w��C���N]�{{�ő3��{\���ĺs+�pg�Y̴ոWW��g�dZ���	%q�dx_�V�/H�L����s�,/��0u����Oe\�۔y�R�f���B,�I�;�m�h{iw����B<���B���5"��՝�9/w51�� 7�?�&�����jW�;_:]�`�8���D� ��B)E9PMi?*XB@��ޫ`^�H�Kn_{�T��~�K}�ș`���]�"���e�*�>G�:Y�W��cd� ���b�_L�Q���_`��#ik�����E2ƹ���#���嶆Q�q�ҩJ�a>���:&P�I��dZ�U;N����>��B���I����k��C�h�=mQ��[�LՋ�V���QT���ECl�3 ��R�^B- �5'��Ϭ�4��8��v�B��Q^ب
�Y <��7�9G��GD-�4�{��+�R�@s�����D�BMi��Q�U#!�ew���
��n�d+^#��A%c@+�V�X����ǩ�;e)(�X^� ���P�5�J��EQ�o�S��E#�Ƌm̉��-���E���҈X��j�3W���|ǁ�H�T��d���vC�-�$�$�x�����;����V����KT����h�.vPWM�ayAY�����v>�+��}�%Q�Wf�,�X�D48���E{P�r(X9��6���Xl���E&��%��	��$��V=��&�0��>k�>�?O��_#B�eͰyF�V,�9����Yx�S��m"�㫮ـؓ��%iP b�BFD��Ĉ�X�ȨMvVdM�v@�x��kR����q��|�z$4�\nb��X�虢š9�����ut�N�ٺa`�o��n�-�8y�4V�[3��{�P�xH��Ǆ~!0{Ў4Pv:��u���6(��:��ZO3:��y����X��mXH�!}��������d�Lw�7��x�E�����K@�)0��/L1~HE�FrM���h�㴬^�B�&�x^�Ku7&A4ꚹz�ο��N���Isf8��~�7����
+�yc=�3��~�l�Q��e@�1=��ڰ?^�Yr&&�*�X�y=5�~yb ���9ʬ'il@A:��p���N��4lF�K�ߵ�����ʳ���%�����?���#;�"��������U��E�4=O�LՀ5��h���{�]������n@�l��~i��>6�}�L���H}��Uu�rGE���+g�/O���8j<_,��O?����׌SF��~��u�OM�Q�O�.hBO�-ۻ��i�����Dނ@����À䝘�T�:l%�0�Φ��Q��j����؟9^=��G<iMB�5wU�p�6[��p�­���sp{��:�}�i�q���NkF�tja+c�a��� 
ʪ��0�;&��ۯ����?Pr.�ia��¡�dk�)�ho^�,�> ���邬%���
o��\M��#~�i����B젬� R��e����QL�o/{D����h��#�U#�eA�I7hk���D����vlj�#�yI�6�������������4Ⅺ�U��Mp�G�wP��x����I�[+V�Wi)#� Z�ۖ�T������27�>�&�	�M��*<��MB,�ʘd���hg����q�8;E����'��dz�q�,`ޙ�ϕyo|uښ���y�M��֨?O�� ����V�(ރx_��fu��JBN1�p}��)�O8���%Q!��j�y0۳Q�O���!gǽ~d�s��g'|W�G�ޠ�$��R���Ĳ���@���wq���̓9H\*D;�L����d"d?*EϠ��'X�k6�`��-k�:����8�0�qQ�D�4���	a�PC�S�7P�!І���P���:
��Q8YJ���M(���XË�@�<::����b}VLo���0z�{<C8�&�OtT	S��G*ٴ�[ߎ��}�^��1������g���!��=�$Zg9��E���;iZ��8�J]+:����}��n�g��W�n��H�d��i���c{�\߳�����a��/%��!<A�dh��ϾG�"#I��z�bvQ�Q0�E���\S��/o��DG�֓q����BKͰ⢔��z�S���αܫX0V|����m�g'H2&F�G]v|[걆��;�����{_F��\`��(N�hfz��>,���u��ЈJ���03�é��y_�pt�ǌށ�aiE0��w�V۳R���f0)��\E>E��w) m?����Y����J�6#�mR8�g]/ZXP����4��Y���jgц]^R�J	�c-��e+2����c�	|��J�Y��sѿ�9���TZ�MT@+2��>4^0�
m��c��I�J\�e��	����14���*w�1:��z������N߈;_�R(�Ʊ\&��T����aU�r�@��G[(c��D6�\tk��,�렅(�D��s^ߐK�;���}d��7�#�,=�-0�i���� �����H�h�^VS��?l@O>0s�B�M����ס�T ��{{!��=�z��o����kXa
��"�%'Ovh�G���F<+�{cK�ջ�/R(;���隐u��~R^eO2c�֕�Ƨ��A༵�8��Ss�a*�p����铵�ǚ����2�S'$,�7#r,I�}h���Y����1]!%����� ��:AFMz���Ya�-֪g=.><CG${�=9�%���"��L��%a��&��y����cGZ
��BG�Û��ā8��Y~t���N�ASyQ�iAS{q���9�?�[�C���"e�Ɩ��j'�ʚ!AfB�aRL���:�%+�I�0���f�|sn$!#A�}9�������%!�fz�\G�Kc&}a.�ņ�"TBr�ه0j�5:��,�4������Ij���E��R��z%�'��
�r ��o�#�ZRBh1{h�1��d��Ŕ�8���;SP���ݝs�R�m\��{O�g��ֽߧ<i�	l�#%04�4�re3�Q[ \膬�2�!��DuX���?�0+~Ϭ�J��v����s^�C�Yl�ug�,�nϖ~�>�7����V�S�R%La�tt/�w���,���1K��pgΝؐU�q5�/�sD���.�_�	�*����ⱻ;�L~_H���q"&i�H#!�X3Ɯ�ɓu��G���ɬ��Z��u�+�pz+��p�@'1H�@�lAv�j,��kPo�HN�&	ɟ���"��ø9O�f>�����{�l׻bGE@jX<F��I!�rѐ�J%�<��~-C�5�Zf�[���a�����7I�?� �p2�s�.-iwW�b�a��
�����c�R��`��T�d���-���	R7��N�5� 7���٢�6����1��p�e��[u=מ*}�0T	��ʚ1��4mD�H�z���}��Y�;堞�F�fo�9�}��1��� ���=,;��e����@�����P'��r���(`��7����z:��e�Vl��^Hw'(�E���p_�k�zO�R�Un4���h���2��*~y��� �'w����!�mC\p�Y�c�/R0�dRߖ���m���í=7.Vd+6�H�p�_�x�M�uA��m!d��t���HH�-�mO(��]�4u�R����}��U�6Z�)��69:H��}�e��������`�Ns�#��H��&jk.�c�*z�R��b�x!$�7�5���<�C
�p����'N���mk���fj��C ��8��%�s^�o��ّ�SC���F#�^����~2��x�������d�MBJ#��$
x靛�5��X!"�n��0���b��_D~ƥ�+7=��7�Aj����u_��E��
��/�<�Xn�}����k=�U����g�E����a��K0��ެqќ�C��������P:��m4��q�����QA���0�m�����T^�P6�y�>��/PsYA��m��>ll�Ġ����w��Z��<A��n��G�q�j<���abS�n�H`�N���(d~?�Ó&�cE8lz��@�[<h\ڣ���<�����i�x@e>Cٽ=�) ��8�ۭ����@{���18%�����x��8b��!�{�L��۪;�;{��nO��'�<���B2�+�f�=��0�*�3�Jj]���"�JHF b���˟n��"��KP�U�6���ֆU��?�����#g�B��Y��
��ĊMVU��
���ڏ�A�y}^�������^19I�W�t����T��eO�5CƖ�r� }�2�d��L?6�p BRķTn�V����:��Y�=�*���[�vӳc�r<�>wP����N�_�Cx�[	�C�P^ƒ���,w;��QK������%�Z�Hbe��i#��{���dyq���� 5���_CS�������M��ޏV8�P�����%{��P]�F����{W!�Ɛ�ya��ŉ�C��q�)�Ι�iZ3k��T6��X�o����!�$�7?3_'U����$�W�Y�F��65D؂�_��d<���ö壨z����{��en�l�����4�$h���Pԡы�t㨚��I�fY\�#v�_���o��W]���u}t@�A�ۗ�A�sB/RrŐ�σ��_��(���;˿p5��y'\��rN�=�$�t_`E�A�v����:�̻%�<+�;-�y_6[\�����J��4$���g	v�;�O����ϙcq�XmZ"��0hg�V�Le�JV�@	E��,�K�Ė�����)x=�E��OC�j�O��{�m�
��@�C��Zz��� 'y��l�m��^2+��+��d�
��&���9��]﮴e����k�d�W�Ro;�/��2�x��u�C#�̊��-��q�ilv~t���P�����έ˦+��v���mHY�w��-���>�a�q�� ^gh#��e�U��ƕ�g�e����п�BxV�@�����i������]�e�(�j��!׬=��9�)EY$p�ڃ�d�h����.���$j���l��6D���O �k:�5ֹ!~�#\����&�ŮOS��/L>��˥l�Z#V�!mZO�U�{���n|`C�����Gq=_��44�f��|�-�Rٳ���:}�E�T��q���$��U�.�4О��%j�Na�0mh�v����K��c�#{!J����.+dJ��(�����s��y��ڤ x�$�.(�u�.c�VHiZ�$���B�6i�U)U[|�ɷ�U:�(�6j��֮t�3�h�Mk/�&����҈��;�I�r�w�j��{\R�����_���� <㋬1�M�.����4L��2��lHQg�j"$��c��i"Њ��+@9Z�ZBH\'[��5�Y��O�_�ŭ2�`��W�'T�z������L,����G�J?���^�3�M���vr�{�<J���-IM�x��.EH��\_\>zs���`��N���(�J�l�4Q1�ƴ���I扮���4=���c����~d�&Fc���X�{���h��]j�`�<kֵ�B�E�Z*��� �4���2��Le�$����nrx+6�G�k}5�=��Cz)��fp@1�ί�y�F�a;'欒V�`����!��K������5U�̉�k3���ʖa'�ީ���6�x�K��X�qN���Pp�Z����X�]����H�&n�.�k��h����v�~����:]ֶ%���2!������|��Q��vX a	Z˷Yȫ�E���N�I(���[=�Z��S�L2��	�^�jpH��bk������'�*j�Yc�%���t/����S=�&���y��܉�o����~�w-�GO�*��Bء�m����/���T�����6��^l(�tv�!��.�~��d#����?c�3�bĕ_)$e�+o����� >�ԕ�Tͺ������חU�p�v��ݘQ"v��7�P9Moz{"� ���=�&�8}��b�,d-��n���"����.�B��5��]�nWe0�-�*�-�T�Y����j�~�8����581_�<oj�`���.C�de~p|p���IR�U�rm�#2��	%�N�p4e�&ZOQ{b�N�щ� @qÒ���95�$��h���J��D��P�|p�(��(`;n� �s�[� �V��}=[�F�r�_���0��kRO�0O{B�m��ޒ�wtPT�S4�����p���UR�E��P&��%������]F� ��?���!���Dg��W�_��c���JmF�Ș͵w� �gj���g�aۨ#���4���l��ǳ���K}�U�D�����U�h�ޚ")	u_-ޓD31�SE���t(Sc!!�; 	,jÏ�2w�q���B���D�0��쒉Qu�凰z�3D҂p�~2"���M$Z@�����FSۄ[
����Ǡ�����a����[:na�=�o�����LYDil��|���ϢT�?���5-'$��/��-���b)ѭ� G@Z�>5<W/��~`<z.�<G"}W�y,�B����S�4ٽ�η�7�U���"S-���gD&�KR�R/R�@U����6���"���w�T��-6"�D�â)� ����M��;v�=�:?D�|䦔i����42��C���G�����%v�WVFӡ������K>����ƫ>����F���qi�z��z�k!f���_��|�ϵ��4E�12���&�<�Z��DH����ޟ�� 9S]�}5�l���l�����@���c4��u�Q�{|s �*q$��~*���\�� ��OPm��ʕLe��r^����@�����?�=���w��D��# ��g]j.��w�f���/Wy݊M�,����7W�?PQ OT�p�J��S��pG��ta_���c<c�̞�V��!	�f3.�@��I|Yt$�U�f;��_[�,�x��G����E}3z�c,p?�2����C5�%-�r2�Ԍ�Jр�vi@�ݯK:.�婢�e���f�>Zut'Q���#��?�_]�;��iʲ���R�q
�GV�B��sA'�-�ǰ5;��M��tɓ7�9m+�鈪��Q
ؾ���q��\)��|͠�jJ���{�?���&g�<�h�EE�������9��_:�.�yٕ���,���:��߉E��i�I%�Ԃy��m��q�kC�~��m�o-`9�-]��È�T1J���+���>6�������יt����%5!)�e޽ 
��d�&;�D^��"ؑ.��]Z�8q�J!z��2}�ܠ��)�i���cq��"�i]W�>�yP"��}o��@��J��]̑�u5	�ÒF:��f��c<�"?,rф�[)��S�D�=��� �AdY|LI���:T4�	Cʞg`�{�vD��w��n��c���2@�����W0%w'��5�m
�&��
O�ùئ�H�I�qj�^W�����W,N�8�A�yO/�� ��G��}�~��#�p1�Rp�jT�߳A������Xg�Wȷ��@ oYTTN�J�HO�Wy�CKj���`�8̊��W	�ׅx�ڀ��w�H��U�,B�'R��8:��n�jE�Fٮ�Nj��fQ��6�OT ���콄!���,�V��.�h���Fi6j���߆CuST$����l�2���5|�Dh�܋EiD�JƏ�#=afA����K��dy����S�* ����ܱ����-~fI���L0�B�%AhV�����YV�֨�q���{e��& ��'rQ�c�(�YP�,�k���Q�5(�����#����\aD��U�9A����8��ڄd0Aڙ���sU��O��(/l&���W_�N/.v��Ja��Vm�z������Q~�gJm/�����ac�:����!)�"/3�VڴJh	;��"�O�r�J����S��;>3"��!r��VN�u��P�U�$��
�U��U9��D���Q;H	�җ�zٔ��׍�,�_n%��[����n1�K�[ >��a���i�/�,�~�l��DP���a���,+e���32�_�f��Aa���Wq��k=����-au����j�K۲�Dn�}IY@��/EO�A�\�R�����m��8�+�ʗ<�+Tx�_F 1D}k[d)g9��Æ�t}Z%W���2��ݎ����{���D��t�t������;ܛ��i3�^��	���:I$�;��/�ǥ���6�X<�i� J�do����o��n�>��.��=��pP��b����S�9��u��J����[�T�+Nk�E��Xvc��6|h&��k%���Q`!���Τ��FG���31."���d�4�"���T	i��xN��!tM(�d�N��գ2�uu�"�5?�Nz�CtT�#�R��o�0?�}^���'��wG�mj��G�`�k�\!s�F�nS�Ss��a��,���P�������FT?�T+ݳx5���Z@[�O���M|bp���fP�㕨���Se�L�B>e%���
���K���d!yk��b�n�l�Y���ݡ��������?�t��>ul=4���r����ܰH�tu�I:�>@�����}o�zI�0�%�)v�WcBfg3��F�~��2d�6�f�\N^�Q&Md"O��Q�Կ�s���{J�sJb�!�dV�Wޔӂ'�XƖ����x��:�8�ğ}���7h���Q:��o?7#�K�^n��#sV`��� �r�z�\�zZ�	X��' TB�^n�J��;�_vh���Jўx�(���N����Bv�8��'�E��O5�B%�G�TnXo3��Jsgu��T%i&uS���+��#��B���G�eu�l"�0T]�]����5Wj���~P,�O�
��}��8���y���uj8�d,js���NP�o�Fbd#��20�)��-B
4'� ��D�R�A)1#�RG[1.!���*V��������EH9?���� M��QZ[';ǔo�2�_���:�kD���@w��m��i�.�h�������a���2�q2�d����U�eٽzW�+�v2�)V֠Y!��ao��C嘹���鏐��K�^[�Ny��ıʎN#���74Q��P%�������>�ix֖O�#;�a���̨m���k��V��v��>��'�!����-$|�+�1�+������|�8Z��L'8s�J��z�aI�"��|�:i<����.+����>��NB8JБh�,`O7��x�NxQ�fF��ѤdDs��^�z�L�a*�JR珉����k�4�R�,=�h�ȑ��җV	E��p�a�C�o�̴_z����Μ�"��*� �����F�2,���L��w��yW�N<��ѷ�j���t<V���Q��n�N��Hy�і��M�������S�̗t/��|Q��p2ԠT� 0��*#����~J����z�P�K%X'���Kʞ1M1sԳ�f���v�$��}^v]QB�<b�1b!�Ĝ��MnNG����c@��
{y`=�Ť��M�'"�]��B>�b�m}g�[>��UF�.{�%�(/+��5S���϶7���4{�3���'|*()�=S6�
��R��Y(���V�N/���|�1��W��n�\)kj�������J4����)�'�yz��u}�5�3 �%��H(#zV*�vu�֡��e��\B���X&�� B�Ծ�I0��{_b�����J��?�M3+�bK��I����d����F��^D%�bU��Ace��`�y�LA^�>N��G,�hEp�T] �ۭ=�Uyù�)}k���+=���EZ��pl�J2	��������MxE��0���:e��9�����z8����&�`��,������q̥�8nU�V���Ȩ�)qg��
�cR�l:�ί�b�Ơ�L4���R����������]��'I��[G0��_����B"���4u�w��իa���ꄀ�wW�2�ԕĄBĤц��)订J����n42
��E�N��+�7����j{�g�9*��W�Cx�US� 	�ɫȠh��I6���s�1t��$�k�^�G�:���8�
|=�:��!��}q�g�J 5��ht�&��N�Vokg^������{8b�+f�h2]���6���������Y��`O�hv��˿k]���������Ee����W�0q���S����a֋P��{>n�j1�c62�3�V�Xh��J���x�+m�'7��!k��@}�;}��U��|���9a�M�5m0��Z������
�G�vt7�u���q�YL�ς50j��_�M:7�W*��3�����8��c��:'s�sɫي����*͵������X<�3.ަG�$���M��6"�I����\"�����ڴ7�su�R)&��2&X����ߴ��0ZC�.i_|��충�xA�`���5��~O�s,`m��Ŧ[���diO�E����<vfD�>��H	/�jDtF9�b�)T�m��B�eԎ�/X=�=2��{���~"֞�}��w�cקpUNb'���"YH�a�Э�����?wb+fBa��ԣ!p��0�^��ȸ����V9�,?߻;�w��%�0z�|�I�f�>v;rO�6�!ߟ��=4S!H�Q+� b=B�ۨ�̷0��]� f��P��xEFAB���G7E#���^=W�8����z���8J_���BA���,�"T��o�_$W@��4��#,C�]���tC@tf�Hv`>b�m�f�eJ���.�G�Xb�Ӌ%4 ��g>m;������Ҹ�*��Y[����@]��^��h�5���.�l#����VZ������4R��q䣰E����L�n.SEȑ��C
��/�/���a�� ��I6�����T@.r��F���`j���:�lg*!�I�,��k
���4��h=��F7����l_ڵ��ra֧�������`̒���w�"%�ȚjU���̽�٬�����AVɴ��e�ޒ^~l~����@׃`��CG~^����!�O[��M<�m�%����9�%�2���{	`�
T�����dQ���PTr�C=T�;�c��ҝ�_��s&)����WL/c��0n+�m�{�Ͳ�c,�2�4��ۚ��jv��Q�rY��a�83+{R��s������'��7ӧ	����q2L �sul��skhDͦ��N hg�#n��ä��GV��rŖ0�o&�BQ_����3�8F�Q�Z��t�D��u&�x��}GQg�3�(Y� ES�JB+i���W����)�N�lf��:���l�u C����A��Y�1Wăؼ�M�Y�<���� Gt�%
0�K�h����:"Â�i��J폮!�9��>�]U)�}�,�:��U\���j4M�W�~�=�c�/�_.�����]��C����5�o��w0���Z.� gLw��`+s� �ݐ�YnMv���a�i�B�^�5%�͇|:7���%ѹ]�����&
j�-��K��n��z�td`�ǾNf��J��?�t�s���7E����5��z�56��}0 ��U�HY���:��7��NU`ln�5�X7��$�p(=e��]Q֒ڻǔ�h6 ��.�n	ۭZ����
����##*���ʅ�����U@8u�`b4{!.�z�G
?�����I�YP��_�c�m��WN�z+��p�����#��d���Q`!�o��o������8r�N�#���!&��\�z(@qiI�E�����sh��;�ߦ)�w  �)6Y�%���_��,�,ɼ H@«ss�A�VK_n
%�o!k ����B~�o�+� 8D�F��-Đ�Om�� g�$�1�#lj09���7$�w�����]�,��$�T���z�r8����e���x�c~���vܫ
�9��E�����qu�&W(1�vx,�A��!C�,W4�b�/D�1;w���@��[L<mkvG��a��/�3��"��G�T��B(�E<������Z<�$q{�A�6��$����QhW�����CY`�|bu;`��h�Du�"u�5q�` L�<A$���3�a�#j��яB�uF�G�x�J6��v�qt�/��e9_[��?��ZC������0�15����K�ה�D ��6>R�	<"����D��g,��Z�I�F+=�/q,�M�zז�i�{������k�L�#�bL*�Ӗv˙d�c�v$\c�N``�YF V�E�{�tp��Y��� 8��?~F��+�J��Ŭ}�O�(J�W���Ūt+*����f�y���r
>��>��nP�7So[I�D�4\��i�2� �wy�O��O����9>��_��u���nt�#�6'w!ce^2NՁ��1���^5(�O��9`m�~����_�����ۣ��)��X�G�#�AZ�kEHG"�=�B.�AS/�����Ѵ���� ��[�M�ud&_Z�����>��{R�]��3Zl(���e��C�k�����A��Hy�;��r�\�E� }u�HoN7\���?*e��'��|����O�.96��u�ݦ��}�j51<���}�
��Bm�O8����d����nY�Z3u�KMbd�������&�=m�K���߻p�� �kX>��E�af�5<�C�\���֩��'�41�O��-#���pDA+�l��N�W���t|�H��0�f,cv�=�K�Da�B*���k�=b�2�'<�����]d�B���# aTV?�I2
(��$\j������9�:�����rWzON�p]Fm!�d�7�{T��,�N f�k�Q�d6��w��z��h{^kB��¼v���>Y6�����^^�-ީ�y�(պ���7���{>��(���zHk�J� ���j�/�` �����U�c;I�� ���X�Yά9��`=�!�	�ub<���:	}�q|�����@��Joz���^�V���#�n�i��a�ӦMt��C�2���'�s����@'���c*��s傰i�t�,�h��X�Q���ŏ���ȯ� �Y���O��v,�N�:�k�'>:¹�6��NH" 5����XR�BX�ؿ�'t^$`
�8Cy����z,_�9�b�=��Q|}޴�/��% P���Ո����*+m�-�}J�?R:�<S���T��n�"'�A!���1V:��x���%�ؿ���y�W�9M���k�|U}�Jڎ[�	�Vb���3O�k����)�X�_�%?�sE��ۂ���|1J2��Q��Q�3hP��y*����t ��gX[�c����3���-��1���s�OGMm��ϣ�S@ 	ͺ��#,Mq�3�c�i�d�� �O�v�3�7����`�MA�M �@kR�7�3oq�QY��Y�t��/Rn_����������]|;��O$n�¹B/n�h�⑟2qF.ƒ\�U1/k�y@���!�uo{����ZU/�~&�/�N:�pGR��!3�D�h��O.wqDggE�k����y�ޑ"ȁ�X��v�}d���]s�D�Y�Yk�^遍�Ƨ�X�P61[�g�j�XX,��p&�`�7`��2�_��A�c��Igt�83��0'J�ߙ��h���Q�%�����\3p��Fg@���fzfS�Za�*퐔��\����Y�5f�4���Q?nQ��0����G��IJ�[�0!R�j�C���jᕻ>�&���"���VqM��f���:~m��{�q��*O9�R�o�>:Y��`��~$���fr��q�7�����h1�>�p�-p���#O������}� �|O� ��6�u� ]��@vrF�NA��W�A��$@v�0�]��I�#%���=u��9P4	wk̋��"���~iGܡz��o�~p(]Q��]1��Y�9�"~]�����Z��`�G���`��[#�ְ?��P0)C��uҼT�N��]D@�{�N�`N����A�~�o �5�f@
|�'���̎g����Fs�5��Y�}!�5Gd~CƧ s;�L�Â� �����l��06�G�uU�U��J�U �����4��J]��6T)������-�iU~b%�0H����n�5����s��u9=6j��[�����!�>|�1����ִ./�tF�U<	���tb�>t*@ ��������#9��i�c\�*A�Tc,с����,W�͏8 S�N8Q(.�'������d
�������|�Bu��W;f�`q�� N��e5��;j�[����������Xxt�y��$��`�0z6�k���"�	s
7��>�#(�La�`���)R�֎��נ���J}�g���#H�P�N��Y�e)�~��UEQny�eN� H�_2�7�ϛ��v(=&��Z��ѠV�g���K#g��5,GB��-ӿ�$�r��-�5D��:�a���:�E�&L$�(ąi����z���>�=�^䋡��r���K���m�߼�2A�cN���X3��J7�{c�*M���1Zd?�Z���tj4!�:��{>q��Ⱶi��n�W]R��ӝ�ڙ�P��x�ν>+k�y�S�`d�{���׹|�H�O��b#H�tI� �U"�Ld�jŲ%�m�=����r�_�����'Q��O�^�Hw�$v;�7��j�jv1���[��];�� ����{�������<�Iz��_�������z��^�Q�>���o� �"�N{�m�$*�_��Kv�줣�ح����\%�]��+l�*S�H�ˇ��E�a�TG�W�
G��jӖ���t��P��'�ѭ�� ^m�8&.8���j�RvZ���SA�T(�-�4����k�W���('~�)�Z���~�d����h8_�/���f�Wl�d���d�i#��V�,}gW0�D#�߽��R�'�����s��[��x?�e/�(���Xf ��3�Q�-/Nv L�G��PZ�[����])�ɦd	3��ã3Y�~m'0P��Ƞ��
x�Xb����T+;_�}Fs��Z�u����.(�7���>AW���:5>�qiD��S����H��w2�	w^x��ͤ,��>`hvڣ�)a����֕gQl��%54�'�7��;o��CF�F�#E�y`'�Q�Chi495�Xd���H0�2 Vg�~_n�W�|k�Yis�r�קr�l�9KW2��2~ß�s��$�7���T ;�9��A*g�j�*v}��T/�| ��!�k���1���WI?A�r��T�����6�?M��qp�����^�0X��h}���w%�)�w��u?�A�χ`��([!��s�Z��§N -�U�H����Z-}?GY�N�T~&5����cѧ���Y��V���o:�����dʞs�D���pJT��Gf^���֓D�x�ƣ7M/f,mP�_]�l��w��g��������ѕ�}�M��}�s?��ZPU�5,��{�h87��-��ғ��=>��[&8�Z��������[���I[�Tb��	󇇄f �;O��,E�1�b3���NRu�*Վ�V�(C����g RM,�����#�苷r�`�xv %N`��J���P�iwN�_��%��+�YD����g|s��$3��}����_���c$@�3�ۡT�p�M�V�����Ϳ++f�@���9|�}dX�Ai����b�'�n���nh	���@h(�M.���q��o�^'�'޵+�/�DX��T�a�����W�9�v/x��r�P��bЂ8F�'OX鬤b�Mx�w��p���$�Y�bW5��sT��F�(����hF=��9��%N�V�)i�J�EbL+A-=3��}o'A����U�wR�8x@���S*�1�K�j� ��!15�I��){���k���Y�U�P�%H�^3�+RSs�}�P�6��A�:�/����T�pN�o�����#Λ_�Q�1����M88>�I8-�&G��-����u\��!����'��H�?W�8��-d8��y>Wt!Ѓ��	B��kJM��M���sJ/�Tf�k�5��4��H�Q�#f�3�5��^�p��7��5��L�\��z��ф��ai��GI3�-���M�2{+����tĎ�ģ䦷;�<,?����3p�|���)P�P��eD�Z��^��%��!A�h��@\�����OL7Ș�;��|� h�r�#<�Ri�y�s�p�ξ/-G��H%E�'��MmR����q���)*��&�gK�l������F�m�f�)��Z?�EE�r����f���u�t��C�w�i���G�a�g��&A
r8�Ӻ���t��nH��Y�̗��!p��nni܌�����դ%;t c<5B��%��k^\{�	�;�����
M���'�׃m��g� ��P���>T���ǎ3��!��� ��0vgﻷU�6
H�OL�5�kd����t��.��oߝ輡�{����?� &�
mv��c!?���:Th�P�dV�n!Q��z'D@�A��ۦU������ϡ�����R���v�?�sN��J�O�7w�gٿ��	�m�����{
�:�ǩm���4]����-��Ƞ@O#u���y���U������(�О�ʳP�I�؁������]�,���l�d��yG[֘����3:b����������Mг���q4�(��}���{2�J�2�?��[iy��K�,_9��_Y�5`i�١�����\���<v�f?c�8#*7���RZ�:�D*Z�����Ŝ�Kz����k�Ot��v��U�2�wt���iV�&�c�N��H��:	{L�A��f?Ԟ�yX�C��_��gUD��'f�r�6Ŋu�<�z ���J��rN�cq���i���Yk�C�y�0�)I����V`8�{R>x�c�t�N�T��Y�i�K࡜�w��L���HqC��N�����	:��z�\�uh��C�4�����˽,q֟�g����l!�f��B�x��I��^P|��v��Ш�(��mIж/��\r�n+a1! �<�MW�ѯ��<h�Z��7�,cR#�R�]� �D�2`��ZH�4�����E��]@.k��^�W�_M�K�XQ��҄l�р��&&	ٯ�ovWr{�M#Z���^���$�o[�W�%���M3ՔZ1�ss�� ����յ�Q�e�r�i]��,@�P\_��R��Fո�=�n�����׮:d�Ё2Y_+A��Hs}�֜ȸ-�rђ�u��������${`�кk���#Nu`�eh�W�hE��g؟m@�1� v[���xV
���)���T�:��];!*;p�qRD�L�fa��5p;�Tj�!�<!�kޕ��߂�O3:긛������٦D$i/�Lu�i�/h��=g�A
���kb�����Чv6�������`h\�C_ݱ������sە��
���uD~R��Jqr�:�P|H`�>1r�:"G����ڋ��R�	�1q��=�b�r׊�Z�g�det�9���I)ͯ������[��ϤR�����!�>'R��^nm�Z,���{�"u>�ڱ�� �>���E��0b�s=F*�=k�x8������o�'A�-χbЦQmn���.����oQVӦ��ZOɂ�l�*�G��it�\����:T�o{W�y:�N�C(!��:�J���d&ɪE�V�L����(���͸���G%�F�ę��'�=�,IE��w�Zf�2�U�{�0I�^��<0z?e'���^~lڙ(�M��";!��j�m����|���s3��pӳ����B�B�`Ks�o�e�_,��{�a���`�Q|=�����&5�5��W�{.N<��F��h������l��&�Uk0�N�:ይ�41���|�꽪�98P��S��_��n�¾��wK�I��Țy�u�
dq]e�r��XɾW�dc7��INK�}ƞ���e@~����Lg����n�����h�4+@C��f,o��z�j���l]�2�\�Tpx�J�#Q�G�n�̍�p���%	L�3�Z���u#��`lM�rx-|P��,�����י�z�*��#�
�׹��2l�Z�m�>P A�Ƌ_�…��к@)��b2���4�����Y�T�=k�t^	c�`>E򮊲�H��YY#�����Һ:]l������ŘNԥne=�4x '���H<)�#�^@~�e7 6�m80ۡ'	V�v��a�<��9�/n|놎Pl��k��N��ϙ�#��c���|@{jrPlcI<��W퉮�
-��P���'�#�����f�P��i�S��#�@cq\�}�L=cɽ��aT3��LMfB�f�?Bc��"��s-�sIK��KK�����W�:����ې��3Xg�C!}��Yϳ;kZ1�,5ƀ�9�f�Mv�+U�?�zv������Ou�a>����%n�11�D{G��n�� i�N_6ϫ�W?�W2�b>��|�=��8�0�:} G�8|k�1��U���q�*�<9�@����&�÷yQlg�����Є�Dt���³v�בN���~&��@�$f�a1��n� ~c����Bq.'��	}j����A�N	7�B��j���X]�!Ю@}�ք�xÁUUC�v2B�1�P���κ9�κ??$�����g!wՖd�P��l4�'{�'S]�wz�6��=A��]X����T4A�<X�+<O~������4I/r���z(Q�]"Q��>�3p�ʖ1��:����[s�y��7h�i0b$�yetyT�a�%4�{�fp*�~�}G�rƳ�j΅�e�3Q�|�)a��*�
��W�΄�Rџ��Q0�$I�� 0�/��eV���bo�n����)�$��C�?9��̀�E�'~����Iy��J�����틪��A2߄��"��-���[�B�Ts*@|p,{3?@�g���O��G۰ Df�:���fh�W *�,m,�N�2c����C���HW�U>��84w�O�������-����ΎG��q���	��4:���Ғ�p��C<�����1�^P+jGdy��+�~-��S��߸ 8��$�WBm�KH�ژ<b�Η|�E� /G�L�ā0��l!������Եp4�҆}"��aG�	ւ�5Ϝ�)<���8
��_κ�3%⦶O���~,!qf����v!�螟�>�U�9K�I�bg�bW%-k�7���?+�a�a\*Z�R��S��j26M�^��#�Ja�ı]����(�=gBc���"����f�v�u"|�0�MFӌ��/�ƙ1S�7����<��>�\�2�+��%�f�A���q��i�g_��*W�;uQ?����@(U�N��[�2��W�᩾�5�H}1ʙ�Î��]�s���޴CX�*�����f0�}HT������*�_YV�|���5��n� ��0���w<�W؜)��#�B22��$���-�j����{>�ͩ���k$(�8jFby��b��h����+Zۆ,��V@����j�)�D�G�|v��Lb��O���%t�k���4⤵�D±7�$ꨠ�Gy��;9Qi\�g�����j��E2;@�:ճN>������v���܉{<����IK��:-g�������Y�҄�u�nS�:�fɘ�Q���^lqf��"P�Ss��I����
�.�(g�{��6B\X�^��1JN�s�S���/�FӬ���7���{�Иݧ)��!��Л�(��j6����m���׽�����0�AA�Q���v%��IǊ��$j4TE���h�<vI���"���n�k�6�>���S0��#Ӥ�Aq+A��%�~o	�S�i�D�C*����Hū�rx9����C�bj��'!ؤ��9˙��1�J�/6T�o>mZ}�%�K�����̀?\YP����{7�f2݈�i�ݣ���w�eJ+��{y��ed��*5������E��c��z;�J��B<�	#��)�qx�����l��Rw�p�[�}����+P�nh��L�>u���#)����m�j�C�I6ҫa�	Q}�qڥ��i�������19Ϗ�p<;�C�o}I"����[���}�pz���x�0<'�yܚ��P�։�?U�0b��QT�Ѹ�e�˲�b
^t�PM� ��Fj�O��b8���qN�003��QB��������:��U<�-�W�QG�(4y��Qt6!�H��zg�^D��
��r�mܮz��KG�y�����/�Ք2h�`���5G=���v|,�u�JU�9��2��c��R�ː�k㪏�����RLu��08�2�KO�J�ز����i�;e���0��K'4�)?+�� �}ϩ�0�TRKί����-ەJ�9�Wp�<\S3�H.���g}c<�O��ڥ)q6O�V9�琸�����j�ߜQ�����XL��&:�;�t���!��VZ4����n�x���7�0C�g�ZێI���Đ)j��+:)*h�XY�k"_[_�����1W�������D4Z���C�eN>��RI������x[��P��Bd��(T���x�&���@%�p�S�n�e}�%����,|��dsgT�X���hޱ���v��Q��c��aAQ���p���k3��ĞXt�^F"���5v~I
u|8��\��N�������:& WO�>���pd?� �8�����	�]o�mU�/��0�'֋��m�[�tN��z0@VK'��=���j��Á���?�{nA�1�Ñ�î	�0��-/M���y�{�t�/����.�+�7���W���=�����d��<*ד-��]�3٢�;ۅ���w��!�?NEvrFޣ��#���~Mqp9����O	��E��?��d��:�2W-6�܁�.�f�ЂD
-F�e��m����0�T���V{��5���W�e��P3X'mӦd	k���?CP�(���2>���[�a�<�.x9Ug�Mg�+z������撘k�<�����QIA�cƩsf��I�X��8I�|�����<oT���oAS\E�j�����~�]Eoc��F�{�
W,Dڟ���$+�!�7�vv��׫o�T��"i�P����.\}L�N��T�~99��m�!�줮�mr!%�@��Y+4\#� q�5���1�`�����'&#��<�)Ҩ�W���%W�L��lb{m,��u���Pr�s�L��N�=�ܺ�2)sۦ�:�uX"��t�C�6BrS�b�-5>Yp��L�]j�����6뀼f�&��\/���y4�\�f�=�şH�%�"�g�� �]�,L���PaRt������\�=d�.��5����qD�~ߛ�����~�$nj��M�E���g�Ó���s	���"�|��W�Z��-��e�p�o��/l}�1񜯦s����i28.��&�ٖ]?�;I����+��J���C��{$�]{W	�]�n�h�"�JH 4��h�b1���w�u"-!�ї��el��j1Y�5G��|0
���9��"��X�;Ŭ	I��y^�Q��e�%�z�m2���m�rU�!B"�m[1����}[A���G�g��3� @&jʋ���PCn��YE���2Nݖ�v�}$��2	6�a�h�s�����R'Esa�F)&��a�9[-���HE��WȮ$����M�<�i+�Di����\�]�'xҩ���3"tS{[�)H��v8��l0YE���� ���SUN������A��
��Q30*Gg��k��{��K?�(Y|ܡ�5����jj>�*��l���Ⱦ.o�Z�c�8��-�;�\��(#�%��"�ϫҝ�φxz�S�X�MS֞�80n�ɽ��%KUe#��Q��Pa�ұ�٧M�����1�z@��.2�y�A,���9�Ǫ݈�z�{ 6Eu䲏��}�v�	W(8��ӡ{�8�w�t9�aE�V�O��p�2� ���Q?`�7��O�
��v�0f
�*0(�g1�{	�H�	jw�n���5����U5��J5���uI'��`*0*����'�1h~�x��f/J�)���Ш���{� �:j�R�	���Zi#2O�j��s�r<��WPɢ�K���)�m����v� �$��p.).�[�&AVv�V}��C����錷w�B�H>3S
��%�ȳ������T���"��\�#8���QEt�|��4`���� �5����}m��W�̏I@m�mBZ�Tĭ��M�S�(@x�.�� �k��k/_ɑ$a�����r��F�}>� :0�f��sЮi*�¬�����ӡ�l�B�>G�brC�eӇ0>;�GM�G�l[���Sg�gTT���N�U�)T#�T\��"4���K�2�����<���MK��r��y!�clT�^���&&�唐��u��R�	ϱ���pl��M�˭�K.���'M��w}�y�t��(�3Ǳ��S�i��S2/2��c���(��?_�C7�D�Q��bT����l�24��Jf��fB�N����!WV�wT�(K�=�~|�{��ڄK���bV�>�E�cϟ�M�Dh������f��0�Cm+�n X6�-D.�o������拏r���k����"7W�t�L����Kb)�DW"��Q�W�W�~"����*�m��8�~Y�^�UK?�m�����ɝ���B��w��ŹŃ�RX�/E�l�iӞLM:�d�1�����6���}����ݐG�nWQM��H6��Y.���"��2c������۪��J��P�-�_�=	@q�S�=EӀ��7�o�Y����#�y`M�^2�4&뎩�IH֢�y�2{^L�����1[���Zd�r{ҁ�,ₕ�����}�A���wƲ2�1�(xб9�Hn?`��F�̑�q��ݾ�*�9J �i� ��"��I+� �yUpْ�G�h�zmG�IQj�^�q\h;�I�]�
�3�_�^�CX���W����UO:j��ؓ1BqzlO�8��ū��`r�����\�S�\C�(�	�d�[��d��X��9f`�];�����^SQ��~�kes=��Q�*n�,��ӵY0n����:�S��Z�.�C���f�W�%'x����=�ʍP�
���u���Y�hs4��.{�\�g}i8�mݑ��l"8fʸ�=����,��?O8^����	�/�D[�lȄ͒B���$f��d֬���]7��-ۉs,��a�Hݦm�5�q�W;���B�bedq�2ѿ��|?v��.�ޔ�M�F�AꨖN�y�E=Ƙ�v���C<f0zyg7{�KȒB@��ta\�Nk�NfA��>q�����G���3�G	�	����("�%���/��nR:fI�7;h/;���� w�.���:�Mq>RJ2m�����&���Hpv��!��?Q��m�1�z�M}��Ѯ0^t\t�N�!q��G\������Mc��CÝ�)��f�s�?C�X�ih��k�{�~R�W��櫋����eqk��@g$8���f�W�{�8���'�]�o���;��^���W����ӵ���ڠӱ���¡�Jn�>�oZ_��:�l�P1w32Cn2�qJ�v���Ǭ�ebA�^��	�F>9MS���OV�m7�ѧ��]#,BbU
C�"��ՎCXJ�n��OlA|���mZ�"΂�za�)Q�e�gS��&$"����oC
���_b	�T==J�Q�����t�0K������b_���;��0�\j���4l�I�`�V����0�Ł�މ~Ҿ��v�Vy�I�=��i�O��[j�2�ڄ�w	�RK���?#��[Βn��z�@1<e��in�t�r&@��8c�����#���r�]jg��+ٲ�����#]m�������&:B�8��"v�ε�uh�6��>�����a��U�,��{�+��>q��h�YQ�|����$|(�4���Ƈ��ĸ�A������(�b9?�Po���b1��g&6�Jh��/��E�=z�ڼ��i/�>�Dt�BT��aq�v�b� ]y���}���ǰj����D���OhOՒcC3#��~o�f���l�Cӭi�Χxy���F��&O;�V&�$�V����.*B-��5����6EnKh�wO,\q".��2U=u�G����p�� ��㝿�Tr��)Нm��fc��V�A# m@���rd�>9\Z�$t���FZ3w�v5�*e����ʝ�S����I�N�;���)|H���W����1y�A^=����7���q��,$$X[֣�t~�� ����٬�k]�������
�:%�%�λ�^�!�Ft"��a�'e�����x��dX��}�	�R�.��b���c���Zfio�Zv O'H4�)F|دW�^�����(�J�u=�2"c��=v���$V��h)��KD]���r:����#otxe΄	-r��s���W_*���`�|}u�e_�G�������;�aMC͐����M�%ۯ�q�WYE���?j~ʴS�il�f��M� �C�X�Z剠���?hWP䌡�� #���b+c1�s}�:��6�YS���4Mt��A��[EQ�5�'�B��ʉ

�m=����4��+9|�<�.���{�:F9d�FSl�^�]��!�C��e��U���͟*��{ذ-�����bx`��;��l-8v�1ﺞ�.����¤��_zl����*�F��6#�O�l������������.k��m���j��w{k7OO��Mz��1m���8}�\�F���	�|���s{��O�˃u�Y�
I�*�Ք	��}6��������^�5鹥5�z��83��D��S��6���et� ��y_ο��*���&%+ �Y-�<���BD�(Vp	�zh�I���F��o�!yRW/R�� Z���ǵ�V`K�ԶZX4�J֡�4^��s6�0���]VU��e�P�L��TwV�K��z��5��adL/���^EU^_��ak�*�$|t��ۊG�5���4�UK�*�W �  �)]���]H�8SN)�J��0uz��1�v7{:��Ϗ����n����Kd�V��]���z��ה3�}��M��h"���h���%��4ɀ����D�F�����b�3���U�ֱ�!fE����q�R�\�-Di�_�����N9X�<>��9ޮT�������1X��:�Ya���	�P���:<xǇ�gJ�����|�pB�,h�0��tDQ� ���X���gyb�"��
��P��(Ͽ�NW���_s3J�َu�z���8��w����#�1��L�Q�!3>ƒC'(�� �}�*�
�v��D�j|������ƅRE�g2	������K�*I����͵{���]����wfI�Ñr��Oꎠ��^���a@��JZ�F��PoF��NX5���e�G�U�z��Ͱ	x]�X�Cp6ܓU
5/~E�U�l�r��P�L`["&]�&���wؒ�f��Ix�9�me�ؿ�'ظ���?lFՆ�f&SS�y��Ih��Y*�������)��%�(����VD�6	���%���nk�Lκ �Jc��la�ƍÿ)ñ���b�R_� �(���)'��Ra���U�+ᕗ�����������9<�2t.u�����;�ӫMJ��VE?����=��e�Yo<� E��C$f7p6B�����ÿ��)D�@uv���|Q�����x=s�����Xr�-�U`�/�g�Gӊ߇f#�0U؍x�O�4��^����c�K��g��m�h�ob�Q��N���k4, �/I}{���Z+T3pU{5(�=���-���Y��u��^%�E����=m���;ݢ��vh���qP"R��b���IʾVj�y��蓨C�a������;7kv���ޅ�	�x���K�/O���v�(��E
.�#����7�����5�
����`�qj5��Rt�!�?�`�ChJ��>��3�#n0PM(����!��/A�=���+GC�B�D�����# �e�������Շ�����7���r՟����F�Z:�%10xf�S�T��I�r�Ȫ�<�S[����׫�[��9z�M��jl�O6��@��akZ 5�}Y	,�A����JO�?��4��̇8�n7�|�o�ɾqS��#]��L�%髿�o1��`�qa5��TN���N������k+��mZ��}�E���B�~�5�Fu0�� �
�EO*dH��߬{^�>�O�^���nc,����b,yBy�L�Gw8bq4��t���%�%�`�}�!],��̽���SIj�s��ֳ��H���]"[���Wo/��#@���ػB���_�m�G!t�t9,k�m�-��-6T����i�Ǿ��=	�<���Hó���k�S�[S)=��0e���M����Hb���X�2`@^�����"��V^1̋3k�y�3:7c(�j
�
9X���=V ?�`cE��3�wɕmk�`���2�{.�?�Id�;P���	FXW��|�^8y��޿:��#�N��Ɯht��͡�2���*�8m!�RSKԠ�t�{��=6G��c4Pb���i�|�G�W?7V����%Nx�^��s�V��)|�����}2��d��[�pr�ql��cM�ޮU�#N�0�����城�7���GQ�/c�
��b����\�?��H	�2�UoZl�,�����F�
峭��[<��c��2�m'�`h޼%E C9ʼTQ��9_{-�r®0��J�.�3�.��o���h���ũ���2�a��-s�(�R�l�=H����ŝ��LC$�^��&��,��e*d*���҉M�S1J�Bʠ���l!�Z����g���j��`]�FQ�l�`����Nv�C�mV�J�_����[枷�ҙ�%hJ)u�pB��M�0�ҵYJ�=�l��7����零�\P��L�Ȱ�Őe+�`$���^*��K��{$�����(�"�h�@Ƥ{֜>�=g��/��2ӱ+��5d��q�_r;H`�z����+~+���J���d��V��O��dn�I|����o��1w,���<�7��s���ZGѦ@��r-f�u78V������s?g�*��L=W}���%�g{,�,�O7Շ��9YI}���Y�l6�(�&r�mWR�	t�	>Q�>�8i&K࿂��H���:�ur�/	\c���Ncf��׮�K�l��9��t�I0^�˹|>E��dzS��6=����BY��9�˽�˿$�}��ɜ��c��ZN��Iq�fyኔ�I�ǤFw���\K�	z�
EG�v�$�WK�u&�N��f1�}�uBIv�>�q��_���q��nGBw>&��L!�|����x�sؑ	M+v�ܕ�t��L ���h�h�
��|_�7|͔�6	��*��u��7v�ɍ���f��>����#�%���^hN��X90��^��]�Y��q��J���QwN��te~�i��	lՁ%����a���?���y!3�%�^-zk���ׄ�#&2	V�P�H
|��T�=3�8 '�|�n�B�X��}Ca�g���ܟ�L�F��['��p+_���u�fn֭�G8���c�Ԭ2�����a���j&R �u�"p��!���S�A�t�y@�߂����}�^:�o��e���2�K���ֻ	���+|}ȉcWzeJj���uhB��0^�۷:gp�f
E飃/����n�E�'h��?������G|=46�YxC��F�VҒ\Jl���8�zbe2���>S�X+��a��mO$�D6��:G�n�	T7��y�-uD��8>X0#��*��O&��!�pŁ�y��7By;�Oܨ�?�#>}���\'�����[-x$M]Y#B#,ޡ�޸�+W�TR& 0�.:��/�[|����\�1r^��q�;�H��";WyE�wo9�a�砠]8:�|}����pA�h��i�'C�k.�{t�	�8J8O�j���էTcD�ĺe�ѣ {<��>�a.��RK�6���M�f}�Q�%�u/.63=D�W�|!'l+y�� ��J�����@��g�k>N��KR�Hކ��]�N	�+m�Dv���p�r�)�����VT�W��
ϼ�m鑼K):�^:�(� <x�%��[q��>?��`۠����F�e{x��h�bOX',9����\�@N%Iv�U^n�f����K�S���tb� :i��������F}��d�:��F���}�����ޛ�b�F �{��S�=,���,P{���*&$�|מ�{�x84����ťI_��uS��Q����|�7}��b�;�B����y�8<��4��������t�a���Q�8���l4ͻ%p 
Ne�s��|���뭒7ւ���0��_����_c��y��C��h�"B�8�̶�m�D�����3R��L%�Ij����P��m����C/��E�4��>��JזJ�0����(�6f��!�[��-��ġ�Ga)�s!���̸c��-��p*��ML�8��HU�O�G�k@wQ%3�����<p�|W�4oT���$�dI^-m76��P6&YZ

8V�La"Lf[�	��{�d�m_��M�q�/5L/ó&��$�0ݓ؊��mee$��P����B;u*¥%{	�eC!PyLW׋{	j̣�|@�=%��=LvP'tQ�Y�w����!�|[�=�ѯ���ł�/�8KۣPǫ�h�`�O,����D��}Ϭn�^��z7��0;����E�p�����4K��J��"%fj��������0��F=��ZW�M��q6�蕡��#�f դ	��������Mq��4����lo}E��\;��gN�B��ଌ�|�N@�2LoLU|w�^���؝��{'�$���Q�Һ���+�
�ڗ���ey�C�s��9��Q`�p���j��Ɵ�*%�?���du�NB���Є�4����_Ӭ6�(�I��G��Wx�=���_�|����(�;L�����{���N�X<=�g�Շ�Uė`��@�o=(�W����uH����h��N^��Kdt�2�:%-����LC���ۭ�I~'���X�aO��E�x���1(pF��%4z�24?��d�}f���w���f-V�Vi�Qh��Cl\���}��6%�����������)*GCi"�}8�7������q����))�`Zh��N����y�5�������_�uW�m���8?�Ȗr��i�I�ː���}b�)8"s��Jа�%NB�z��Ag�5��|�7,���2���w�3Rn^ƪ
�S��-t�v2]��H]!�c��`���D�l�p������a�r���6��*Zn}�n2�Z����omC�8&�("���0�(ʕ��0�G�X�c�U�-���(�N�̱s	8�*�� ��tj��UuM�@ߩ�A����]���M�aC�evL��3e��}Yd�L��'�$�hܹD�+G��-��p�z���!�p4n��CJ�!���W!Qr]s�].5�[ꂢN~#2�b�����jۓ���M���f����Џfx)�47�(~JM�W]�w���h+ټF%.�Hs#�!Y
;Ґ�,(�L7��f�b}D�~����4278^�����r�GRU��`��n ](I����M]E�X�3y�{����y�f��^P.�K���Ȗ�����g�
�h�
�U��G+�ũ&�\��\�GRc惏���XA�,�3�DՃ|�IS�$ �o��A��F��r��7��t|q�π�M���c����/�)D�I)��V� �*쓉��6���2`M�;�a5D �&;+�'1��q��V�~���C�2�\i�ܔ��7��L7)HTxe�/���!\�t,�*8gx�C��N��q~�����=`M���9�7���1|����?���\r}�:
\�
��B������Δ��`�: +sd�pP��D&�h�<8��d�����C���PmG��y7tX�um�����Q�nl�e�$��	P�-ø߷Gȳm��7���Bb���V@�L��}������%%.$  MN�&8Fu)��9^hk��8	q7nizq��X2*�_+�o�t5�)��i/�ƀS��CM����^��Ya�*����;a�����%sK.���7SA&����n&\7��C	��F�-Gs ��c�3���?�
�,�:���]}\�Lib�2i��m���$�p~��`���l�UZFRC�� ���]D�(z�z�I�m�I�\�	��c�y<�Ρ����ɧubr-Q�g~DZ�%Y�NF���8X���d��	B�M�l���DLD�N��Ɛ���-���ױcKU����!�/1FIR�7!�7{#�uXz�ݸ�0!�\YiuC�C^>�`u��I�ș��t�TH�����~��k`1�r 	�=ލR�2�I��u�4&�n�9@�\����� ym���O�rv�!����~����_cwg��b����������r*�Ep�����p�	ȩ]�|$?�3��~w4�sf�7p浿��y���Q�D�w\�sf��|�w� t�8�<�HJ��0Vj�9M�+\���sbz]`5�:���eU�6�qf��ބ@ܖ]���D�Lo���d�|9(2��� �$!b�����B���T?c¨��D�#��VTO�����M��� aMG/��L?��>��,�b���#�6A�F���8s_ ��_cl���� �`}��9?X.��,fͥ7�V�\OXlOA�[�c_Էz#�}R�]k�f�5��V)GDO��g�[�e��*��9"���t�k�
v٤Ћ�|Ϋu��)����z2u�,v_��e�~A�_������Z)�*L�QU��Lg ��|��!l�#�jh�/�r;,H9���A�����%��}Kْ�:� Dt�K�q�^���>=�Ȏn���a�]�|���N�9~����/���U)���b[WZ��	~�H�@�)Yf7��X?T�Ȳ;��U�!t�fvM ��7y]���j��p��<��z%��X�ǯ���l�e�% >�\;\ǡ*z�<�S��X\�iW.��؎Y+_��y�������Sc�����󓓰5��|D��E��t�i�xZQ0dV��P�9l*��p�vd�C�%|"���!�/���N�:yH��7�rE�n��2Y�,z�Ό���훦�ٜ�H��j��qe�
v»�6�T2;_�_oP�a튀��5;�8��{O|M"PU&�%�y	�tO����Z�ᙝ~����;�Fz�?HvK�i�����w^�tӬ�	�/�L�q���V��PS�%��>�)�MhAb7Tw���&d�qP5�,l�����ɿ�Z( J��pM�?�W�����m3%X�_��`~�F)����[[������.% �3d�e�,L�����s�w��GC�q�;E�t��l�ep��V&Mg� t��	��TN}$���5���9>�o��U"�O�Y�Pt;���*�-�� �H�y�'mӵ镽���H#��i ���y>ZOkb&y����D��A���A�A�+mѳ���7s�*�1�PLH�O�����C�O��:X+!��7��#n�'�ĉ��)�����A[ϧ�\�X���X.e���	XA4�GME�8Q'O��Tt�;_���f~�>kڏ+�z�Xi�\	�����h��6Y���`Je��^ZL1�JH�J�lH|�	"��{�^�q�>[�g�7a*��a$��hu�eH��_��N}=�:<A�����qر��WQ֗�5`��׌z��ӰD�P�#uJ����z���j.\j�Yi���<�~v�@��_�b$uT�D��;��S��X�Rh�/HU�XY'�f��O6��S�?�(�'��%颒�u�%���z�@�_�#�o	��f���n��9���
ɱ٥	�H��Go��v�ma�&GR�HQvK�F�Buf
Mp�3X//2L��,��c*���v���q�K"k�E͑M.�۽��&[T�\UL'A+Z$���l��j�&��:e
�'Yڟ�g���wl����)q�(^_�|�m��EL�xOl)��&�q�3����7&C�.�kN�m
�	j�]�i�A���.�Ъ��yЈy�:�?���g�j�~@ ���Kl��x��"sUMc ���3�=�B$�bŘct'��GG@r����|tP��C/=�ڱ�{K�G���	N[xQL��P�b^_ ��nS��U���>��gC�K43@����/랯���)WA����Ѧg�'��r��-�X)\�Gj�(�/.���
D6df, ˬ��>)��	� ����*`l�a�;=�w��@̳et�ƀ�cU�78h�Z���'iVD�GUt�[�4�z���a�3��W;�Q`�K
@����L�_�P"�سMIH����CN}��>��$9���b��F�lo��Kfۍ��"�"52���"Ol������A�J��.�#z�~���=�zؗi��߰ן��2������O��H�Y�_�vN�a�ΞF�-��-Ϫ�(:y$����+FG�p ��Q�*�.(O]�̬"�Uk���2�olE��+��Ѹ���P]�l�~jr�JE�5|W��6Ns�Z�����������b��}��f7�� ���&��m�N���`�t��C�mZ��m�C������\�?K:OPzE��\d�(AH;"aҵ��'T���y�%��N�����.��I�_��� �2�f��YQUK�hfYV��~�z�%>�'�	�S/&�Y�F�8��fd��ąZN�<�T@�r��f=q,Hco��cs���v{5������9R�ڠf�i�S ��"Na��}��J��x�� ���B ��83DTx�zڻ��8wm���+��~��SԨ�`�e"��G����h�XyN�>��Tr,���ef^>V���5���(X&4��D�]|�Xm�����XT�N���@rB�rwJ]��({>�L�|<g��d�x���^��"�S�P���4���}��.��pL"��u� vi�
�k����ľ+j�q��넸���b)	��?���S��O���/��$��^K-=�������� }�����_;��q+-���Ms|�B  :]n�F]{�������Z��j��t�-�ޢV
,����$���D;@z�.�@��c��{��1�;-f2�Vm�`�`����Q����!�%�⳩�f�'�ņ��l� L,��#��pVY�x�/�=����w�����c��|jqv�� �
�����Բ.�� ���ڛ�g򬙴�;(��0�ʿ�t^����K)>��Y,+��xнPi�0��.��4���b�����-�X����,���3���#��JI�Q�I���V�Ygz�N�����|ը���|�E�р�.o�\�*�E�����py'��A �#�h��Ú��7tz�T�*�A����Hx���oX�O����k�#��#�0�m]�Y�� $/��]�.xEc��a���橰6?�n�#��?�A���Qx;0��kz�J̵�J9\�&�G	S>�b�#���1��&��}J�^7��lֲ�]�OH��%��I�}C�
���m���9W�7ǵy�7$Tm�1}��@�� �V�=zx4��
�;3B��)V��?�W�;���N�:8���c���׎r��T�M�UЅ�X�4�Y��`ʶ�B�D�ږsɲq�j���A����
��E39��]�T!�:8C���_O,[o���>��Pk���������t�s��y[1�^^;�������p+e���P{���o������de�E�1�KMg�e����<�|Q�1�E����Dz��L_���G�@^��Ʉ%�׾�w��֖�X�"�g����1[�$�W�f�-7H�3+�p�	�}�@V���s�s�
f�щ�Fa,�[�m�|ho�u�v���6H�:�"�&d��Y誀�ືU\�|�P���&��ϓF��lr+�����R&־�)%�Qn��_�`>f8��$���\��˔����v	�p"�_M�D:��p���ui�YD͈	P�$
e�:��xN���|�%�S�zl��Ma��ʿ)O����u�w ����Ȫ�$OB��TÒ���/�������� v��-3J�ܵ]�İϬxY�_�����b�$*�98Y�z�8&�M-Q��FoHN����Ht�;�מ��
��Uj�u�^�y��T���Y�4�K�U��M�[�u�<2y:G���i�\Y�=J��ʅ�� �*6�����c���q�n^'ֵ�pC���~���&%Y+�L��"��[V�"�Q�ˎ�ͧ�Q����ׂx��@���F9����t�`�<Ո��INKǽ���ܮQ�d�P5�u�䋿��P3�0	_��懙�������P�"������!�\��O~�q+� �����������ߞ�Pa#F��e�F���#��YrWh���&*�K�L� Z�����a��T�.��3�d8_�b�<�I4�fsJ챶��,8��i��{�v�����I��LMs+��w�}<	���6ݻ|R-k�s���U(]���o��3���[�>�+?ޙl�7E���Ckɖ�X�D~�F)Χ�t�s�	�|&c�����G�H',�X�8o�	�L:Y�]^QW��L���Q�Wc*�Ħ���D����)8�_a�p�\n��&�W���O���<e���U]����^(ހ:N�Z=Z�$ub��"4u~8��%�����ڬd�?`Y����(���S������A!0V�|�S���+��m�u�v?�	@�0�6��mϜ~|�i��h����<�4�Q��"�$[M�I�`���"=R��3H1� ���6���E�)U[�,��/�)���ϹYpɀZ��o��3�K�K��
�q���R�o�R��_!̷�7GFv92�,�[۶��%Pߗq�Bt;�~S ��q:�4,MNm��(F�X�BR#����-�\Q'i�'�.Y���a�#I�q���lơz�u�Y� ���i�~�7y_||Ύ��q��⥫�#,D_x!#r9_?9���=�W�\���|�;�A�&�ؼ��o�PY��3��Vf݉�����m���a�w����i	��Еʐ���R=1C�l0�@²�rœM.��.�HV�hAI����5v8i*�.��|� ��y�g�1C ���f�RL�5\i(��g&����ǘX4P}�p�a���C��B!�\�|j}�Y������.��1t�����6P�ӂK����Uh��`Y U�
 V��*��]$2$�����6*˓t,W��Ī 'l~h"On�<���۲��9��?#Jg�c&��.������`7������f���Q=۫�(�2�������&�
I;�T#|sПj�I��d�����X"��!���hԙ����Lk���\��M�B��7^1j�^%7?=vB�ʸE"3��9�bl걟u�;
\UͯJ(S8g+#P�+�_�%�̀�P`v����C�h,ȸ'�B���i���%6�aj?\ᾄV|EǤi���� �;�PHL����c�0��4^PS
�Ԑ�*?�)E'������LVFh���}m�!���)�o�X�w&�R�E)�,��Βݫ�[�<׸+JIwfy�MsI��o�ɔ��k���k�U�@ַ�T:�ʲn��}�ˬN����),�u�/m*n�V������>�9���sx5��*�Xի!J�欲4v��7�Oݎ��0������ӹh�HM8�����J<; �9
I:9�{o�ff<�h��ݿ��U�l�K�g����zԤ�&��%ҍ�ӝB�lP.���� �bclNVڏ2�L)��ֿC��{NkY�U��O�L샌���L:W� x�b�⚀w �TKȜ�N�͋6҆�:�~���//c�vA,���y�=�/���؄n����#�t�Ų{X�Z�O{���4�>�R8O_�L&�aE_�qcSس/j�d'�M�T��]v[aoc��Q�41����܆��@1R�Q#ǂ:k49ߎ�6g��P��qPk�Cd����~Ssl˒,�'t�5�ڌj��f��EY�T:u��J�#X�Ƣ{��=��;�ŬֳBg�������9�߼xp�1��WB����j���D*<����@���־�B����H=������1��s�T�����Wz �� �.��kVP(�$A~[S���d �(e�<����ǧr���?PvS1\: Wj���u�"�6��ƻ3cz̯��3 ��ӝ��- ���ض.?#�����oA�{j���&�����}�e)Cڴ���L��K��fv�J���S����ƺ|�h�\��'A���O�L�5�����ߓ�kI�s��ӹ�W�ܟ�q��d��Q{�^�r����-GH=s��9fQ�Un���0�*ţoU�NA]m�YK�d��`6�`R��.bz�y��%�We!RI8� 8`]�u��kx%L?�Z�Gac>�+�>F����\�o�ZѨ�&����J�D2���g,�H�%rq�7`��%�gT4A��w�S�of�n�� �������|��r�������K�p���&���헙6�>ɣf�C���?�\�V�G�9�W��V��г?�jxs5.E�@G8�ð��Q�6�np���:s��G?4͉d,�Ҧ��ɺ�H���U%��M�7����0`7A)��*[Q�trh�B��P��D���ޤ̑L��6�0G�$Ok�\o�:s(�]OA$��K�YJA���:�Z0��S`45���O-$�{�EI��Oxc%>�J���q�Z�$<j��S��@%;��\&��Ն^v �9|��	�;�	ѾJ��(�є����,ї�ˁ�!m��	4�R�f�R��7I���M{�z]����1�!%rg���W:z�5w블H�A�N�;�ἴM�EGq�Rq8��m(����&����P$Y���N)���+%���D���V�����kI�/�v�`Z��^��ӈ�Q��k��0RS��I��*�X)���,n�"�\L�ѥ�/���KG�����Z�ڀ����w�xa6�V3/�p�v+ ��j�O�}���J������]@��Ɉ�,��	����(E���WЁ-��D'Yd��v��a���0)Y��0Em�3E�c�kN�ߘ�C�շ��-������,*�����p�D�Ζʼ�X�w��E��B;I�[㡶
*��S�|R�����.��V�$i����6��7����1���ز/�-�oQ�5��]�X<���%Kf')l�Y��tW��^�9���9~;T�<�)�) O��W}t��`�!
�5�R�i�:{]�u�?�_��rm�י�lnJz�l�^	�m�Z.��X��M�y��J!s�>3 ����B[��e	@o%1v��ׇW�QEy�5>W���:&N���Ȋ�{"Ձkr�!fv�Z���s�@=_A�2͒c�����2�[��;M�t��9(�o���ޗ$<�z<6�w<q��[�D��V"�R x⯭������ [kB��r5=B)ڡ+X����s���-���s�_ V msnk{�D��~ܤ]U�3|��f�U�y�ee������V�.No�3S�	��%>SZ�vS�փ�6�n9| ~���j6�95j2���j5y��;W�Kl��ؘBz��=2F�{�����1��X�6�&�mnP����C�����t�r���/��M���׫W9u������ ��	}ޗia�:8�����(�J��v�����=�sO���#U?��1�D���s`5F �7yX��v?u#i�dr�W��T}fj� �Xw]�)Ѱς�0<�c1�T����J�����*G �p�|�Ŕ�TK�`���ŝ_�R>H+O;?B�mc*����YV��eW�zWB�`�eKD��~��(��c�-������\=Ik�ʄ�����\ugcI�a�d�a�uT���xL�s_��7u�MNL�*�݂�珍>�`E��l�	�Si�(�!	��?�|������L�:�f�#�y}�������J�"vl>q"��� ��d�Š��H<Ζ���˶�E�,7�o'f�>�,̰L�қ`mJ���I��$lQ�"�C֫օ'�cU�����%��g�XN����_��M���`�Yk�&ь�Y�i�S�CPVOΊ�w��N�4�NC�'�]7��gE��`�`�-l��\U�x�0h�����B,)��Q�VK��T:n��i4�� r�*�f�V�6r��_����lh`��2� L��v_������y5 ���/�_�Ƿ��,+*��z���;����Ͻ�
�(�ֆ������Ѯ��=����5|
���u����2X|;<����RR�^.�1�DԊ�UZmg�k�Ѷ�_���$#��i��hHqg\n��~����$�|���y{/YJ{ozߣc��}�F��j�?k��h��w��I-.��;�m��W��3Xͷ�l��F��xe���h��c|l!�OuH��Ҁp)��O5��4n;��`m�|����A��[m�u���i��h�3g�����|PV�
q��>2�t�W�~0��|��<�x���ɐןa�E�N�(ծ�i� P��T�Ox�忯mgI�`d�=ļ��T���i1�]�6 ���<M����b���M�>R�!�3�C�',�0,����"��Zy/���T1�H�� r�%��@5�zC��^�a��5�$$o����R�/fӑF�ЌvW����jɼ'����w?�ϴ��	�u�)'�����1����Ȫ3E_�[�o�S؉/Ԧf�?���4;�{\��t�����^qQ�6jb�����׹ڊ�i:�С�<�%%�dpj���/�ض`I7�w�
q�>���`
:Sp'K����}�������}�����BRϮ��΀���B�7CH�=�y~�N&X�����j �xl�����]�z$~���K-��^��������V�+Q�aD�Q��%3೟V�އF4f\�>�W�i1��W�b����m����̃"�M3Uj��2��P������c�����Q�暇���D�-�?�>y�����Q$�n��j�
NN������~����~��~�'��}M�V	��`�m-]�4��EV#-�nG��6�~C�x��n>������z��c��V����̄����B�B�fك��������V��.6�e j�s��A���Gr���T��A�B���+lJ��l-`���%�ɧ�?/�|tex��|3{#5 ���˛������	k�(�!(G�<��q����>�����n*��kPoo#V�c�F��I�ŇP�R� ��Dg��wD��Sظ�����;��,oIz��`��N�hۙ���L)�9���Tc
xzZ9�����V�l8	�
h������s�j(?%�G5��=_r柺�}I�$�2ݮ�o��������(gD*�Lv�r庩�ėd$�A�q���I$���>:�6Aώ��y��/���e�����?����{"w�N`�S�$�97�$�_rA�u5���n�����3�u�(�P��z>P��f��y�����rkX���} "nSB��P_�ǥ�~����*}p� ���
�z�������_�h�m>�4�P���I.�u�s��c�'&�!d�[�1��?��U�H�R�R���"`d8[���6�N(i��vnf\bz��(&z��YnQ!�-Ð0�T*��fľ^�\L[�J% ��\H�&�S�~
&J�9���xHJ�y�H��B����2<�w�f�(� �ER4c�U��J�r�l*Tx.p�$�j�a���;�B0���6�t2X=ӣ�IH��K�Y����-����7�����q�� 0�b��ߍJ؉��G��aC	{��	��_Y��j�Z�e��,#3�{�q��~s����?�i�6_�(,,�>��N(D(��R<hh3�ә��:Q�baE¼
N�u �x��x��� �n�Vp#�����N'���姹XM��Z�i]�Ǒ�Ԣ�,�'|:��(S~���У3��*r5w=�����ʖ��;~�z��ENش�W��e�|8m�����fcyh�4�e͍���!]4�sd:ק<��<H�,�Hԕ���H	����Ec�������\��+�1@Gj�iR���_������I���ʘ���N)��I�������Η�����-f��S(_�y��	��o�L��8ӫ�GD�%���
�SK�Z��%c�B�����lv��>Y����S�z����¡~�s־��bo� �6�]M��~�͢����E�op�,s�}��:d��sO�r��/���΢VNd�̍��Х>�`�J},��;�� +��T��]�p�#�tIhn�ol�ȓ�� &��=��@p�iD�$-pɲ<�L�J��+��������}�*h�x�����-C��l~v��c$;f�M�|ޫ�Z��+�z������L�砍��v�w���z\3y
�J�;(�,�����q:�� ψt-b� =T@�@��;�����8�����K�)��Ntl�|��]���"u�����qyӊ�Qe�/fd>/��g��nmde�-�)�r^�\�lr �3����=�K{#�g�;j�1�^{�蝊�.�h  �i�'�-���-��]���l��{�|  �����ф7�W?J���f�۪�=��li%�~v�4i�Ap�+�b-�f0(�jO��<[����c�Ryi�a�ݞ4#�^
�5K��t
�s/+~&��s�����2�t+�Z	�z~��?�DC�%H�?AT�+O�_�D��M;;������~����J�vS�����浙�#�*���������e��'i¸�J� ��B��2_�uT��h�^�>b��R�A��)7'�������!�n�웵��8�v����F�%��k�gcP(��KS��K�j-��w�z95�4���nȀ��0�m��%��!����#���^#�=e -cޮɪ�z��iQ>�?�f���mꂣ�m5=������
��̀G�9�5�ohsH�guJ�9L�fM���y|ߴ����漢�[Co�6h���P����_e�p>�������f8�xXMM=
�QO����IAT��r�5>�.�.x\{��9	����D�7��-3,���83�o	as��	�=�:����E� ��㼗��inJgL�*�� �9[�׳�b������Bj^���0�N�K���Y�a���#ڪ���w�I/B����Ĥ'x�}�G��{���,�9}��Yy�9l��Cb������{?S��k�w��	3�SI�����D����,�~M��1Sa�������U������E����iXᦰ��[˃�MG���!U�eaٶ������M�LD��4����Zq��_�%^�I���q��b	E��	��@"�[ſ+(�(�3�[l���g��)�1�TL�I-��zDF�I�n�B��������!Y9�Z�Sğ6L)թI��A%F�C
j�C�U������#yeu��rہ��:="r U=eȼ;9�z )C�46�ǆ!�h�M�7g���Ȁ���	|�w�Pl�7���|)�[��Gxp�i:L��s�d��Z\jh���~O�!J?�q)��"�i@n�t��{MdA�z��'�G��Z��cB`i�p̍��:%��l�=A)Yv��s"�X]��?H�+��u0!Qɻ�����A냘!s����B�|A��g)ɃEj�����vE�-���d�h4&n=��o7�$��ǯr��
�`�'_�!�Z���6�<���Հs���E�����)��c���*$0.�
Ziy�R���=+�F�?��?�T�.WJ��h�]�ax�6qg�[,�6� �W���	���u�N�,M|���
t��OLC��d�d�,�J۱cSc�D���μ\���x���}���'��8��Q$�S0�ĳݵSR?ĥ)w�(��o�〰~I;����ŗ)a�jx��0�~�pA��c��<`S�t��3��"W�����!�Y��{��\��%��x$ů~V���J��EJ^!7�<w3�h`!O���-����[�����Oa��7U޼���(g��̙?��lQ�m|��G�	�����n-ulu�B��028g��i��{�z�5k��2�C�%���ǔ�;�f[��.l�'�ʃ������盻jR�����]�\Z�gROS�w�H����dg�܁̇<j�!X�/����ʪ2M��dqi����SZ)��uF��R�րn��_%�}h���p�������j�̨.�I����Rw�P��ЎT�;3���1>����D�7\LٱXN�UV�S�,
	7Ho-�UtJMYS����q�F�Ɯ�����ҡȵ.M׬ɗ�&���q��@��;�)� �NQ��䢸wB!��c�cw�P*�����2�7�8�*P�	�[*lZ-�y-Im�FA������W����RP�x@ά'뽮�p4%z1oT�.E������$XO��7n�RU:��Ф'/��Q�S2��X{�N����c0�bM�6Э���o8摇'Q��)A4���\l�)����r�s)0�e~*��zm��k}.�E{+�NiTg*��_�)�߁RE{�?�}aA,�<�aY��S>>JŔY���� [ʀ���ae@jO;0����M�R(�q@�A�7���6���ȷz5��}��Ϻ�W8/R*�~���t_&bҪ���&�D�m}����o�5��y\�<�����"�/w�Ia+���>8�[��)ڻ�?W���lT!�1��9���Ji?&�7����6al*i��M���|��V�O��W���ĕ��@�t�;��d�tXHe��|K��XB��L[I#�W~�R4?9W<ⴛ���\J���/>��(�#�=n��;,3fשˈS�76�I���r�;�7~�+����תm��P����('�`��xC!Ʊ%�J��e���9^�i�<ڻd+Go�A�(*b��h���x�`VX��a�K[����+�vֵJ1��2�ıP�
��`u?M^���C�dO�,�Jm�zy�ZL�����6����O⾿m;�AB��8���Mew�r�bȀR�egr�����{[Ai��8�m6�L
��6l�NMb�����r��?�~��_�G5�9��"qV�p�r��D�Ƃ��qF�y:��]'X���ϯz��Mˆ�K88�=`�&Y��)����:���3"c�B	�ｧ�q`�^d�����E�=�a�:aRK%04����Q\w*�N�����N�I��cKj�r��H���ZAU����Rz@�����F�+��f��O0�T�kd�=�B��S�f'9�rn~����AU�U��5�#��o����&m�C�|TN�"��pyA��_�����_>��k�	9�h��>=���-��1�� �S�[�6\N�r�����]��s�(���y�P-#rm<���T|b�F���E"��)������Ikc'^�8Rh%������h�K�,���p�wj^� 	�;H/0���P����]Lt��u��ֺ�S}.�<:�Z���Мn���eҽ'g�x�6���]k�:�^z�/R��6{K�*V7��fj�D��Ơ�Ϝ���+_�}�VX�b�0���t,�GIR�Sn�5�(�ON?rj�dY���x2>Va^�^NH�9�|%lu-�'b��^8��dD�|.�$ZPS����&�W!W�aT�Ѹ�&!W���� �:��R���u��T%r\�[��q�Xkm��9����A���jP�=uC�U����Z�-�ņ,\%�����v�T���Vj%���*�E��;rf!���/,A�6}kC�?,��̗
wר���$��3�nv�߷C7�AE<��q��>�݊N����5
K����B	��{��mZ�4�s�i�G(�����H����j a�XNUR�U �\Îu�~�֦c2S�ˇ�lT��iYb|�9X�$����}hA)?�a����~�%5�<����G�n��o4q�$5���QE�Q��߷ŖElI��x�'*%l��u�<�U���Z~HGn���&F�\ɽ�
h}���U8�|a{��c`-ot�=�l�����5!3�jO�\�7՜�?�z�Α"�ըR�zu�Ռ��g�z������"L�S���]�Ϻ��k�ڒlX�8�����Pr��XD��T�Г�d$��C�k#+Ợ��.= <).�OJ�2k�Kb�sI]���5����@p�ToX��������[B�Ҥ���M���s�骰�E���~݇H��#��>�K��{`dlksg�C��9�'��
�-ős�gE�|)`��'�z��7�!�¤-k�"ư�DNu}��"֑�g'^Q��6?���� u��u�v0��(5���	�h]��n�13�3�9=��v�s3O�����zR�����&?�?g��z\�c�b�+��%Di���ȍ������u*Ett4�Pkx��M01_�����֗���`S���CG�(�0Cǎr�_�RPʦ�MD_5����3�R��
;��:*+_L���a>�`�t�7(�rN�l��/�Q�P�]d�=�;�KNl�(���w�k�����\p¢�\XH�͂�x����u6C�^v0Ȥ��Y����<C�#�e�GA����@&�W�|�a�%��@����{�4�B�v���2�nO�"���:ǘ�[\o�v��5���@� �M��k��4:���j�r��v%��$���K ����*�a��I���T�l������/�.#��������JRh��`��E�����!c����ҋ��G̊g��](WwR���=X?�@����u������cM��9#����GaS�E�%.�	ƔÄ'��+b���d�����!ﲽ ��sP3�Gots���c}"t+g|"S�G�@���"�օ*�]�5q��l'"g�W�Y���#���pl=|�0���sbz$2��qd[���Y	iG-�$ _ք[���،Q	�P�Ȅ`&Z6A�M=�#�K޴�SӸ�r�L�F�c�N6K7�C?�K�x��`a4�1�A�H��\�����������W�Y�@�$��1����Q3��D }����Zͷ�� %�BWX�0���,B"�ոJds�f�"g`��lџ���$p(V~���2H..�@�-��s��EQHc�[#
�[���������L���|jq$�^Qkx���V.�����Aڷ�$�u�D��Ka�T~�dCiT[�S��7J���[�`�?	<��>Kd���ܡ���q@��������`�δ�k�6�)�%U�7�ƗͿ��c0��['F�X�p)��c!�G`aA���]g'�Ci��i�۞��9o���逻o�� 6ɬ��lc�<'���F��&�Cn��o)QU�ζ�C�fX.m���@�
�� ��8���eK��g�n�Hω��B���T`�Y�Ӛ��Eu���Db(�&�P�2��+�̪g�7wz��?#A��Z��j����7r��jf�d��5a<��R�@ �<�K��@�.�]��`���OȬ�z��u3��Meb��n_<�*jn�'?l�m������GX�/�˟�gQ�ڄ�yM)6�m�i2�է��tϻk}���͔;�,�5/V�W�A&����)���
$<��hp�`P@�ҟW�TA����@�O��T�y���8��#�1��y����O}DE��j&�L�Dh�K���a"�Z{AG�/lh [��oK�Y��)��:+��V��wc�9+ݭ�͐
���e��%�V��G.�l}x�E�a���J�&$��;BC�2����/j��K-�S�s:B;��K��k�zA����g"#.�$����ȍ���l��9.p��]P��o`c�$�vUKؼO-���Y�/wO.���p��\;�w�z,����k�\=����Q�,��ŷ	u�|�I	�'��Xy��z�ֵ�����+Al������2�P�u-[�|��/59�ˎ����BY�W�n��ç���0�@�R8爠��NUz�u&=�w���>���;�dƴ�ɤ�3���7�	ڻ���5"�x�B�u*�#���M���:��σ�
���{T�ș�R�%�%�E�U���|��oW)�K�����p�!_8	A<Pi�O[|)�
şg�ʠ��T�9ˣ�e�^s܊(q�XmY�
��L��K�ɇ�ƚF��X V��"��$7�b�ה���ogp����8�D�����B6v.�dJ��D}s�~K�`����ՠ_Ջ2�\�8�~����Xxp�e�!�&�#G?|^Vd@�L`�/q=�2��E�d-���!F
o}��4�wk`Q��W1cl�`W��qpUy��!��aL��%���$�����Q�%�4�V��#��9��I1^�(�49	�ח&�j�z����ܸ[C!ꤎ��T�"�fӶ�¾���!�#�F"R��f�ܨ9R�D�P������uC�L��V���}�<�q�Q���X~"�}bZ��)F�EȢ�6��~��lm��G�������`�0���Ēm���LӮ0u����d�UA0{��5K��:�쪯�,Lj�=�i� ATGk���/s�?���:�Ɓ�n*�����tO���7�a�8D�>N<~��
B�����FUSЁ�դt��2LȲ�Zh�<It���:Sg�R�A�T�?i�i��}�
�
�q��i����:���e �����t	�<5�S�U�tRU@�n��YGB��aR#�wF�@'H���EJlR�]�u)7��UoX�Mc��v�K�u����k�'�9�4��������x��dڷ��>RбQ;�H���;��G�@����k2]0D]~&O�Uꀮ���QH(��cJ�
���k�SM���r >��/.FF�s��{9��<�1	zM��vu�� 5��`�YA�����<��/MwG#�k���Uw����Dm-	A=p=_]Ϙ�����*�5wl؍�LO"u�2�� ������2Ô���A�WV�"W��`H�uq#�hU�.*P��[f��Di�N�7%�&2�`���1�_��P�@8%�Q��*	+��lD��ӾO��=�P�/�ܒ,��T�W;b:���<���B��>ߵ��Մ�3�m��;�F�sk�#s��$n���O�?� ��6��ѿ�!_�m��[hS�o���*L����oP��h/1��[���%�+m|Q>�z��<$�g~F��Z�[�z+�X̝V����T��Y#8n��	��0�g6�*�#KƦ��1BFoC�� ��!���L�??!�s����w�K�לgl��5|�G+��b�*Bi-�t,��l�c̜p"�$�b@B��G~�������Uv�(؜��w�a�ŝ�o��'��@k������GOX�i�X�Hӕf�� ר�����{�hvQWӗ9�%ɸ���Yh���9ኾ�P|&��� tֲ��X���=���=S�싁�q�5�����D����n��G�g^d�0,���gL6�C��tIW���N������u�3�E��3?�-vp�3�l���t@UP���P��T�@�_�^�!�c�x@v ��ߠRyɀ�������&(��ϭs�,� ;L�Xw���c"���k���ӌ �qg�H�U%n��<�u�=yd�_9������^�g��d�ρ�W{�/ ��}o�Hx�}�y/8p>�	d��Tz�ֻ)v����˪����Ha݃"_��V��0?>��7$x�L(?ֆ8�FXL��?\�p{�Cc�e�M8=�����GB���x�b�V���������PIi3��n��إ�½����Xh ʩN	�����Y��-�(�cq�j�*�D�+�+�LT�E�q:��9 �t�#ȹAѰ��D�yDu��W��gm�"H`^�����J?g��#K~l�V;�0�U���!痪�:��(D�Ǯ)��0ڤ7�K�z�Pm�=��>�=���|PL��w}m�x�x�E�s$?A
#w��K1�keL}a*���*�V��]'����"m��[P�yGH��߄%;�2X���� \1���X�N��A�e:x�x``�Bu�m�������)�h��ew�ڦ��X��j�J|-�w�Zv�ٙ�a��'6���Keӫ��o�����0H�1���!5E���/�$��4W�JVi�3�;ݟ���R�p�RI��!˂�ɟ���V٘ӽӂ�͆�Bq�dk�����_��W6c����r����e�f�W�C���ZA0O�*�q�[�rj���)o�1&Ɣ\��5sG�%k�.[Ԃ���Ṏ.>� HҴ��,@��U�5���}Ƞ�B^0bX9j��,`��~�l؊�'�n�J˰Yb��Y���ж��Zwf2�&أ��3�ڵ���9���CV�늋��=/5�5��Ɋ	m�T7�S�7e��ʚ�ͱ�.W��Ѽ�vĮ��^�����S"�Q��ej�r��*�fV��#��f�?oV;@�T1܄�v��>����/��L5)��zZ���h4s�.
��NC<���hK����V1�Ers�lbm~�C�a�J�G@�y#_�'GJ'���L2�� b'�2�94$�-k����/;+8�Z!S5���@��(�O����jr�q�\s�A�[6�<���6HW�����'(��[��?��X����}�(�����{;�'v֢a�sD��9.�$�q-���Z�<XV��釻���W����@�ak�hp6t@�6Mt�u����f#���1����%�S}ܾ��=�h����"�b#��N���]A:=P�l��$�υڳ.��I'ޥ�����A��Ft�3¹0��ѓ:�|�D�8-;��M�ua�6�;�W�!�n|d�$g��a�n�V��I�j���C�i��\G,(���y����8��8Gk�{����Ob���V\�W�	�$�E����D����ȵ#��o��T���'T��'���o�rW )TᑉO������R��
�������/j%��5���Р���?K�X�e����*�L��T?��źX�a�V�����ʎ�(��x�{[��N �ל2�I���up�<?��2y�A�@k�,���!����̚Qi]�`]���Q��!4�4���[˻L}\�b���`φ�zu}�,"O�Qʌx�0��L)�*���ah!aW�^�ױYd�ֹ}k5�Ǡ���93}~�Y0B<O�I1e���_���D�V='D��_�����]&����;�v��b,x�گ��J����G��|��
�2x�z��>�d�U9ڜ7F� .�'�{��Qg��Q3�l����T�###%��:nh��&ã���uM_�%�ŉF����)�bU��?u'����������͐��������re���c>���T:Ã ���e�1�D�i���^ 8��h�j�6	{c���� ��3Ɉb���8]����h��9�VB'
���(���WƮ��0��Q��"&XUC��p�B��s���;��=L�N>3�[�bbe2M0��[Z�[.���a)�g/��h�Z/��Ѡ7宁F�T��w�U>���U��c�ݢ�)̇�^�]���Rxp����bA)A�9�m�Lg����"�������gXf���kG����Uϕ��k����\y&�X�XU+؎tI0�\�Dʙ�9!յ��-d�wU��S���l�dQO�\�vitd�.�������"3k��]=�1
�5L���cAC��|��_�@\!���ͮ���ت�l�Ƈ?�.l#p�7���;u01j*��Ԟ��<?*��=a2�J�M��i�ƙ�Ԟ'v�.�S�6[נ�u�E:.X*��6�����=S��oYhߦ,f�h9��zl ނ��Bk�ϒk?c�\P�e�r�q��"+���e֩I3N�[��� ��TP��ք����(?�w�}y�:�1��/��N�� #�u��Px�ݐx�s�U�P@�m�L�Eh#�����I�X��1�}��v���,sԐ��n�O-�NO� �R9R�\I�_��i��I/=�A�����F���ۀtU��*0f�4))��V��w$��M��Ga_���S��שkÊ�`����?B7V�i2�^�"��Y��@�����|�j(W㤅���bF��9������!$������Ś��lW�QŪ�Q,�}9x*�k�]iI1�%�|���L�iGVf#|�x�L����B�R�;`Ļdg�8q������q�10S�\��ɭ>tfş���-|���f�	Y��[����%�g���
Mc��;N-	P ����K_���p_>]ͼG�yjB��
���F�e�ZL-���ř�+K�$Ź}Hg������<鏡d����� o�Fڳq]^ {��\b���B�4�F����)B����R��aT���)n��+��V�8�'}R�ut�
��Z�"��������G�"�A�	�h�$ x׏�d
	˾x�FG���u'3jF/��s���^ G�r��v�����]��IƘ�T�z��7Ptx�#+�G�����;�Dծ��&�N=�Z�j�R�휊��j��t�)e��cV�e��9^H&튖����jǽ�g�|HPnj�߉��6���Sж���a(���揉�Y�U���˭��_����d���be��u�r����O���߄>��W �li�jP�y��о刂������M�;����ٿ ��3(�FX-������j��?�Ei��i,&�$�f,�1y	T1�1���L�40�Ї���Ta���4|�������(�H��'��9����������d e���"�^�)1�G3S4��K�_�����G�{�@{�y�I��>�M��v��ؤ��sX�B�-��Gm�>��e���;�SB��U��S-�Z����v�-��]L>LQшӽ�Y���<��>� �=M#ޢH�H_����'��sA�십�?Im^���^V��z�l9,T�b1�,�5
�۩�����S�x{�'%��w����o�%{��·ީ�F���:KN�^�q+!$s���I�ҕb���3!u����1���Z���i�ŴF�"�Oǵ�I�p��(5if�(�.w��(�mhjW_IAP'j��}ʧ�o���I c˜��D��{� ��:1����q
Sw��-�Z���Tdu�Nf ��^�~�Q��y]smqrX�QB�t㨼�F]MQT�4�nX\ꛥ��B���w��u�5��]kG�����N�/ �C�mi���˭Ct`t[_;����~���h�񉝟�E�u>^����/��[�����*�I���=�5b֒�mu#�.��DA���6�EU�G�ว�=����/&A[ I��Oc��.��c�zq���)T��ύJf� �e[��_�Y�����������D�G�ogjn��v2��^��C�2���G{���g�2naQ�6�&�*<&%h���Q���uK�dS����1����;8��;PN%a����m��S�
I<���DO��QT�G�*�;��Ko�wS0�O󷀭q��3��f��~�2���n�B�/2����N�i9�Ώ��v+ӳrՉ��r%���B��w�j�ܕ�мZG�O{T�� FP�!�WG`g�H�8$|Vh:r0�k0��Ə�U���(	j�-��[�,��DT��2�����������Q��?�����7Xb��^�ǰ��?�~偺�`1n�f����o�- ެc�3�m�]Ts�^F� ���)��~,�?�N�J���RZ��Ȼ��-yUj,��˿�+��(>x���.n���w�1�z
Pߣh��j����r�Ql�}ƾ�9� �)<[������l>�:;�<P�(N�<3�x����|�0�[�FWW�Ж��#�G̪�����3W���[�]����F��V3�^�O��N��R tu�^#�|J�~9���[I���9���p�dP?����c�/� �����a=��g7��dM]<V�O��%u;�$�i!<}3_�x�!C�ۧ
���T��)ʟ�D��m�;��d����4!�|k��iQ\��+\�WeH!���f��(GS-a�h�r�],q�w��|�����ER	j��8�L;���40]p�<�أQ���5���h��(�j<ul�zN��1U|�� ,'J��b����J�z)�Ml������)�`H/����7��j����)���dح���I��W8u�?^�=�MH�.�)��BĄ@�4j\����Cy�h]7���'A�XQ��Jm��i�=��L�N�������~��8�B���^mHw0ğ��$1+c���b�6�7��������PGc<6��mܕQ������B$*~?�w&/�Z��dP�D�Wy%[M4Eh�}�Q��H�Ú��b��WE�E?��m!����$h�j���Mt5Vո���/dܶ��)�w�_?S�Uv�%��Ȫ��\IN3C�Q�T`��-nbr^kfy=����Kc�'��AP[AI�^	W���������?�������vz�~'v6y�×�sW
R����;U�.���qR;��c�fU�,u���?� $��+��]q�9��/�D�	Y�[��J��*�����*_r���}��@{�K\*��z�:�����z���9go�R���y���_�7e	�'���}�I��G��~��y�O.J� (4��j�u{Q�O�%��G�~�?{� %�׬]��0���%AF/�9��B�F��cFj���7{��j*��e	�TŲL�a0#O%�@as�6��i�!��dD�)hҼ��caL�Bo�QS�Q���x���d1�ۉQfO�էm�m���x�k���M�j�]ǌWg#%)�(+s43Đk�b��1��Kh�������ȻBq��
��(�p��N�� �}"j�(n��fL ��|�x	�\@���ԣJ�Y9S\�J- ���,X� �9�����~�e�J�ۯ3M~�G��YJ�i�;��ܼ���>-c�זF�H�|6�~l��v���,��HKY�,P�i������D�pG�FHw�P11���= ����n�Wղ�h/�jOf�U�R�<�'���m�d��t�;,���N��&wE>Yh�WsP	G-��å��?v�ԲRu�i93�h3T�:ũ 3pC��5RGnP��D�ZfJ��T���b�W��}oε�9�F>Uĝ����<�&�Vg�@�)����Log����Z�2!��h�5d�]�ޔ��.�������HU�*��[<�v�C�ǔ��j�' �L�����S��جd���Jko\"P�:��C�=e�q��*�B�UE��&�~v�ea
��搰��;px� 
�z�P� ��q����G8\���!<�%N*e.�=�TD�m%F�`b��j���ۦ��	?�k�6��>�MTPxv��el����Ku�0�u���"GB=Zz�����.b4��*�����&���ڬ̡vhP���E������<p�DF�y���E֤����d~�y�I7�������_��^EM� b��09�G�#*����/�'�5����B��LP��������M#V]�b]~NƬ�׬���<|}����ҵ�� ��[?���iE���ɩ��������+���s 3Q
���Д�THu!��xbf�(i�I����6#��Ͷ+WM2��VxS8���[Al ���B/ɍ0Mq0S�n2mb�ζ-x�}���s*�ɋ\�r)�Q��gӺ"�����F��A񍹆<<������{�Ϙ�
H��0���E!�W$9�B[���"��[�; ��h�o�Y3�i�O��Do�.�5k���R>\�K3	x(ʓ�v�!�� �_S��G��@s��j��ܳ��&t�`�kb�A��1�`�}��#��T�d~:}+H�jH�<��ic�QD�#���|R�#X�bH`�����N�9��Q1��5i�.�z(��B2CjW�B�8���Y��7񶯢��]��\�rvP=�CT4�'=e&Q�t�?[�1����!��9��M��,�:������M7����k����(s�t%�ڛm>�6tMԻ֍�R$}�TÛRC��z�F�U�����Br�,�:\��go/��|��2�YdH-�GC�5n�,{�O�Zq�檛# �N��N�i��D{u'�8Z����J����5(���	�P%>�x|r�\����a����׉խ���\V��:Ϻ�X��!����o�x7���~��Kze��6�%�xH�W�����BZݑI�ZX�`�yL�S����$�o�&�	�_�*bc�(sO�D&�
��O�����h�����dJ�\آl��?�K�G�5=���i�T�fI1)$��l$��(�̯���l���Q�1ŉm� Y8h��: �jn뼖p�$[��åC�N!`4WD�1��F��)p����v���ڔt��VeeEb��.�n���*A�2O�R�d�����S:�_U4d~��x�_��Cv�%�V�$=wG6�QcU�k��#;2�$��"���Gk�V`���9ǲ�䏃�l%V]X�<��-��+ʤ�m�K�}(C1��;|\l  ��^?R�wom��A͈&�0�hw[S_�|6x-Aa	��h:� ��g�6[��������oq�kXI ͓��v�`K*"�_�B��F�y�VC�u��9l�f%8 i!�|F9KaP��G��B>��S�$X%�I����o 3zBN!�Jg�u��G�%J��jb�a݈�0����-��r�b*ϫa�GE�<��>2��x ة��1d��S/Y��@A_�-��E`��b��_�G�Մ)�w帮�ӌ�Q��N	W�GN;˥�2��Ԡw�M�l�D�K#؞al��ֆ�>�.F�)�@R&d��-��F�?�N�X�p�`*'���b��t8�l��/��;�`� �N�$y.R�u��W�ht�Y���� 
;��޷�?�7�x�D��`����Dޜ?�������
�؄�w�SQLy���ِ{����'�e=o�5�&|�Ǽ���7ם������'��F�m�
*�5�6���r����'���Y2��i:Ԥ�7�S��zh���|<�+��̃/O_���pD�Q��ƣ�j�g�Xߧ��M����M�L�)2��X��:����Į���c;�ne@�O��*MKYءV��5%-d=3=lI���ڳ�i�����q���*\���HVz�Z����M"��ɹ�E�ZF�f�Yg*�F���<T6��	�0T��/���=Ax+�q��@����V��$
ޅJ�� >�y��M�i����S�!Mu_Up�r,ۏD級���63�Q�:+M��vw�7�	Lq�H������r&��tp��]��^ڸ�S�_�s|w��p�K�w�Ww`����2P=I�ދ�HZ��
e���Q�Cyk{X�V��&�g;	<xS��z�ا�b)����t��X�$I��"൶�﹘ �_�Z ��ɏ��1���0�_[�k��Sw�[Rq��7I�?�kk'{<�
Z8Ф| Tb��\;�A �9�rv��bs�m(��ڎ�c�!*��T�dqO�L=����]��L�D��a��W�T�v�E ��W�g��#>ED��дo�%v��ICU:y�2��Xq�������Q�J��D���>ɥ�$�ʁ�`8���k=QEIdʽr>6��aDe���n���=VZ�]����P��(�􀋛�^��������uc���(��+�O�팷��VC%^'��v{�^��K��7��k��H���;�@�����X�:����CW�B�Cf�O����݉-�{�Å���y���W��E�R� xh����4U����d��]H����YL!3��69_���w�w�E��cva
����I<;*�Y����I������( 4qa��eQ��TG�C0i�X��:�D�6W8�4B�P|TXi�C�7fa�ш���`����NZ�ޣy�4i�������|�׫�J^	s��Cd)f�7V�����z�,P�sʫwW�|�o�oi���`��/8W;�P��a�䳫��(��؝T�J6��'4������I|c0R}[�!r0�m��d��8����%�Z
氦��XR�٩P�>`�/�z�����n�NنE�+��m��:Z�G�W����9#6��R��r�}�M����&w�HF_�9�#��vDj���M;��aQ����'�,P@l�B�oÞ�c3��3;���4��lQ�Bf���%���*�V�n��&m�G���5U�@�d&�������KX�=W�0"� +��Py���`���5�Zk���)��7�AU��|+:�aǽ����|@�3SP#�r��M��C�1�'5ϜO��K�� 1��k�í�K��z�㛶��xtַ� ����<����b��־����ʇ=�"dȒnO���V�߰!���FF����cB��ͣ30Vz�[L����[i�����s
������f��C�éG��L���fR@��*������0����:X�Y��B}��m��Q��7W�Ǥ׀�c��ŜWZfR(�7�hT���[ 0v�Ń����z��g��V�a-��=`�0"��4 ��ڬSm�#�:�{\��V5���B\�F&�}x�^P�-
�nE)㠍&�KnT7j~���P��VM\�ȍY��x��.�1�H�=�����N~�L�qj(����^t�xx_8�.��fH��#j�
��d�Ci'����*��ow��H5k_�kq�L��blr���������Ky��ӓ�����&�FM"���%y�j��$1�χeh��an�x�<p��`��kk'"�`޺��̻�3���L���^��"�ν�<����D�j���Ѣ�ѫ���E�/;�'-��J��օ/`�_��^(���o��,>�R���;߄ �������WJ7����e's�s\���Kc���ރ�'��^M��m@��H�ą���	*�A*4p ��`I���W]ﺫ��{:��7}�dھ쨨ʯU��Mᅪvh�-2�+�Mￇ�,A���/���)+3ҽ��\&�S�_f����"��k�jv",���յf�y���z�=H�3�@��k�wzW!'7ڴ|��$:&���ڧ=΅ʐ��:/^G[.�\��]]��,������Q6� �˓~����V \�᧑l�]i��o<�p�'���I���|�+��7�~f��͂�S)����"�����`>}����QP��\��E�{.[K_���ZM���h
�k��	ϼ���_�Q��[��RDj�H�bl�*!]O����ձ�G#J =b:`Қy�h�jS�3MWYit ]k���-c�R{�N��\3�5���d=^5�>���>��=Q\�?�:�=��1(�:{���/�,`�$Ѽ��1c���a3ծb>�w�iE�`������*��H�Z�p������}�F`rA�j��Ý�	v
i��{�����׬��=j���b_�l�\�.O��*Gk���z��9 ó[���僦���@L*�8#�z��g@W<���L�.ˌVí��K���
�B�����I.	c{�W��*>В���9`��S�"Q���y�~��3zvY�9����/�v�?�|"6<H�N�T�K�#�ZK.�Lk�Q`Zx�½����}Zk�}A��Fr�P��|fG�aɥ�O�e�����#�x⿩��NVLṧG��	a���vWp��o��*�s�L�ХF�	��7�4�h� .<p��3�ʩ�6��K_��ͩ�ML��Fj,F��]��Le������d�]��@(��~31Ĳ�8�L$�@vQ	�<k�N�5J�9Qr9U`2�t�	���偙���x��:�����T"���C�cFAS�4�W�ָ��8��?)w�m7�A�/T�ҐTZ�&�c�At��46���u�D��V�ɻD���"w+s�R����[��� �"B�'NR^>��ee���%����"��e��$��k���b2�`���]��E'2��}Oz�]��Os��mpӺ��Rٺ
�3�2�����zSXکݤ�׊S�)�SCݣ��W"�')ȱ�&�xJ��c!�b�S`/ ,���02!�t��
����<��$b?Q�<�n:�?��}i���!!�gM��g��F�u��a`a`�Y�$��I����m������U��6\p��p哹ʆ���X�����W��2x��;^��W� !+���j$��������c�9<�'(2.Px�Rtc	yآ�r?�i/iY�s%G�"���������:�m�΂/t8�@�<j�1�UH���L�;;m2���>E��{��7�����}�0����p�H#�����h��:1��%�F#T��̞�L=vTL�Wqi���-u��_��s؈���m�B2	��[s�~t/���PS.z���{���R�F��Y�;��&�q+���ㅣI�}�C��� ��4b5�8v���<�uޕ�K����A�uەT՞As��ݼ;��	3��R���|��Cu&{ !��Uz�Y�f��_�E�uy|\4dū,��sթX� Cl&vP;:��󥎴<W�`���EN���CNl�x��AheOT�G���߲�+���M�c�9Q�C��@��A�_��T�c	;�c]?�ܝJ*�v�]\ͳx�d�0��z�=����@#�(<��O��4O� ڊ�����0�#%�b���\�hM��K�?3H�Wʢ�)t�+
��y8�s}� ��'�_�$����oT,�U�(@�z_u�5�k;�M����= ��,#�ܷz�Y)C��Xtrݒ^��v�K����M�u��ͱ���m~%Z�͢_��_I��D2��7�m:�dy�}g��W(��# �F1�낎�����R�o��s&��-a�y����}N&�̀����2���/����]O��Hw=xo<w9ҵ6�4�Y���#� �Ġz��x�VQ��!�A���Po�1��_{����i4E"ݬ�{�v6|��`[`���z�6���cX{K��q54<s�ޯ��2g�-ٱ�����u��i�}a���ĩx(���74ݼ�oӇ���SO�VMm�����gW�uW,+5V1�ZԈhu���񭙍0}�.�׵[Y��W�\X~Z�P�w'M�2��Q�J[%���n�����8�L���z��F�j�u;> �c��r�w����!C�.��&�+��AC���?��k�+��W4}� x�Ie��Sy֠G�*,T���E�1�����'C7ЉM}�#�&'�[!�GQ'�=��%�D��Y.J�(�$(IDg��-�*�-��X$m�
,�֙aé����$�if�)n���g���q�v��m��&tc�s�T��͖5�� H��D��W.:�a"ֵo2�i�'܂��b�M$������Gv����I.���v����ڪ����Y������ti���?ּ��}$n7A2���S��H���A��ᯫ��@�) ��eSՌ�1+��x�1q�q5� U"C/�����*VBߨ�j�~�O~(���A$H��!קfB�|�1\���P����ď��Zlr�f��2��O�t�c]9�ȴ�љr��&hy��f���m��6&�0:fO���}�)�؆<{9����t�XVv��ľy���l3�5b�xFC���WѦ�7h%��i�o=��(X��]!Z�K�2S~�'O�å�M�O=�3H+N5���siI���͇�Mt��-+9U�9w�3��!;փj�2�����W���S���L����D��j��m�����d�5��'��S�$켜e���Z��5kA�ʻ�N��0(-UX���V�}ѝK$�}�\͐I_���{�Ϙ!����J���0�v���,c��E���:F��F�ԣ�>2l�"[�	�6�{�GbO�B��>E�lNN\���Bl���M��P�ϓ�V�����q�)�%��GpU�'�^D��d,$'
N@R��;�����������&�w����z�[ H�a!�T��������_��Q��d��T�=�0Zf@�1�AZX�&�f�%G"o6eɝ�j]��9�ߎ�&Q�oI�D�y���c�A�S���"I�Ѓj�[���y�$�Y��G O���;�`@*��5Zu����(������*����)��h��\LOS��<�ږ��w��u����2�����Q.�����<���c����Ȼ��������,41ַ�N�K����!��q$1`��>�������x�<���U�N3+��ھ���К9�λJ��HMm�^����D;�BH�w�Х����g��Q�в�]�1�^~�U�om�r�_���z�<�XFR[���������=���C�B[I�EN?_��m��K���3��:�@�4�Ȩ�.uL�{Q��璫`�(ܧ�>����\�W�5.���s�p^#~dk�*��g.^��p��+���`Y��u��ni�Oj��`ߦ�:�+SI� �p�Ӹ�^�%\�w�V(������[�=��.'yem?�G�e���[sw��Ӝ�[�d��wo�v(L_�o�#���~�ϝ����=�䡝C8 ίe�Ư�yvSS[��0����Λ
�v��EBL?�j�vd��w��V�S��5�P�=f��	Iq��߫�Q�#����n{�P�����0<��9�X�L�/{�n��X�VH����ؑ%B��+A�^��.����_ޗ`jx/��?�-A�I�]n,�&��ہ�M��*�VS���/:z � �6��G�_yfUQ������+z�C��>��������$ ��c݈�HߨE�D��}���dLTjS�,�+%
bVχ����D��	������[,�Z;[�҈]s��5pp�THRf)F��z��C�7��A\K[22���y:�'_K��/�b�ڑ�*eQ3`v���~�Y��M��k�7Yk3p57џ)�#y�c|�f!�^���r?'�)rdQ`��"؍���*R����6��4-��,+c
0@1��{,O����8}��g�2Q
�>�a����x�hp���o�Ȧl.a�`^�T�NjV�1^�
8�X�n�c��,hd/�.���u��Õy��_�Ƽ�]6Tľ�H�N�#[�Q��R���������"�΃s~�=��q܍u�%T7���n����h[
_�'��� 'a�-%.\3���fu�w�O`bw�b�����ط0:<�N�"������_5w��'��{��m�e�"����;ԁA-?�^���1���ĺ	=i,ݘ��:�6�'�c\z�E1$�c5k���]��Ӳ�&�\�1����$2,�U3�d�ґ��sb ソ^�6L:D`�m5�c�u<���ŀ��`�����ۆ�B�G�S�ഌ�K���8��U���]��	���V0Tk9�VpN-��lT�z'�vJ�d�S�E��G-E�^��N�a��3�Q�.�q��pf�s�&�ZR�u�XW�8��`����i�S���`��R� t�r�=N�<o���:���W1A"��f~���K�©�l�FE�\�p�Z6�����k!ΗHB52z������uT�w�W���dP���>l
A � h_I<]"��\d���tV�-��f�S93~	?��YqC�V����\��"/�~4AqS-���5��W�$AKl�g!�H"^��,BW[A6��ލU�T���tj}���+��$�.1��� ��u��X��ٔ~����!h])���C{�?(
���_Ρ�ك�'Cy�΢J�ŏ�(~�	�V�O���E�r
�-XT-?-���v��z�E��f��i�۱�y*N����w�����]%0�r��	�Y~��W�}�~�q}X�6�?|ɜ"�>��{B�j̉j{�V/��,T��dL\䖖�ݞ�x�#V��p��N��v>�|�|:��/.7��g���Zs=
w8t�{�������u#$|�¡b7��Fy��3W@GJ<H_�`��f�1
m]�}*}-���vV�M�c��l�<�����b�F��Y�
���Xz�ĵ�~��C׈�j��j~�a���>4�����F�"|���n�Y���l�9�ГS��|K|�j�b7�%G������d)z�h����W?���"��,�Q�T�Ȋw5|^��p��u�n��6Z�R�ꛡ��L�^�6OrT��!����p�~sV��~��C��Eۖ���Je��b�2��#��ʒԲ�Eyd�iu3�t��5�&��e3G����G�G����yCI ��j��`�6��E�ҧ�j!@?}�1R�Q��X@e��BT(�I���W0Q)H]���X��E_%g���#�E����i�M��=Wɱ���K_�{_yG%�a5��G(� d5�����ϕd�dN�`z";��܈�x�$5��rQ��K{��/^{�ɩ��e3��5m�̦�����S![gᗿ�m*����I�\1I��~�z�T��N��R8�B�skM�ֶ�	�	�Q�Hp&|Eʬf,��L��X�P��`Q �,u��}�)��P^��b�D��V׾�dW�PGU�C��*Z�K>�(��du�Mf`��]���s�^�Ê���36�	 ��Ѵ� ��߭z��DЀҴO5�x�DJl��%�2��
g��6�"�]�VD��`F��+	 C+�h�ǣc�>g���ho7��3Ƃ���i/�>��C��'�7ɷ�YS@�Ox�m T�Ҵވ��qr��9�sV�O���06��ZF�"ǒ��p}Ά��Rd(���bJ�%���.��e̹kΪr�-�󕡻�w���U⌄돝I��N�]��h�;��T����y	�h	ӷ+9�a�rM��c��W0!9ا��/���d��߯.��e��b�N�Z�/&#��҅��;JC_cOf9�\w�1F��M��mI�o�M�}CJ��/�KO�r���vX�[�j��=�>����i�UJ� �Ms�8���"�+Ń�ԪEX/�y!�c�4
����bPvw�2.2E��һ��$�uH�I BX%Uo;�=��XH�/>;�V7�*�Sc� �|驆��Y��X"��U����m/e�v5J���A��~=���7���^��9o��=K]���5l��V�R�7�1F�ȼ�Y�g�m!���dޏJ6e�F7��@����dA��=��x��Њ��ͷ�����1���Ќ��m�l�������3�[�1*�����(5*��w˂xGˁb�#� �n�{���v�H���R�@}<>%�6f=��w&  t2���zm��%�1�[b��V ,%�@�M�T�?	b��qF׃.�T��;�-Q��}�>_��CR�e��q3��h���l�+��̤����9��1�B�:\-��4ӈ�Q���=�ƌ�,JH�u�w��6�,���z�i�FV��SJ�ڛ"�vh�͕��`}��O
��[��؍}_�3 d��� � Q����"ӱ)�w���[�{ �F_-w�=��$�n�"��(N�R�9�bs��q��7�-��kN�Y�������_V��0�($حQ:�ش*�&�r�w����W�ع�!�jg�3�K1E�}��n33SZrl2Z &���US��!"�>HA�ˉ"ٵ��@R_^(^*�Q�H~l���{/D������V�+�
����39$ͭ�� ��o��ı�����s"3�f=�f}5e}��<��5K��i|��i��aAc�@;�e���0t2e�3��=7��r��md���V6���uB$��7�|���xj[Y��B�շ�:N�;�l�ܻ�RA�����m�CU䥗��o29!���ڏ�e
�^i��)������<�k��/	��W_9>~1P�W2�d�r�Y�djM���jߙ�#�X락��e�0�d%�	]wB�N�[��֫��Ǭ��?K#[nd}Ͳ�Gr�`UIO}���a��G�����kKu^f�9�=ԻA�G�D�\���\�)��,������]HXr�r�T��FZd�c�8�"Ѧ%|�A���+��ȡ�J��o�P&ϒX��`C��M��!������ܘ���-�b��ܦ�<���3@�-IUJ�_h���1yF�X�]�^ǔ�`��M}��'�X���DvN,���|��[�}f�t�1�8>�
2���h��%I��M�!���оb���Jೈ�bD���s攒KLù^�%NLڻ�V[�]��Ȳ�@l��]��F�Q���*$�~F�D��&��/�i�t�w.��Җ�ny8�C;���Ҩ��&ȡ�O�v�K��s�z��3�!3&��5}?J�^{8�.?'��Wi8�Jm�����֤e^)�7[�n���*�/��y�W�L��{2ýx��p�ְ�N�m�-O��,\���Diz�m��]#��z|
�*�8�(�E�s]�2�ŘU5��N�J�>y��(W♼Y�*�0S;G���SaOn�o�d5?��� '���9vƍ��,�R��n�-tȶ��$�
~^��Ri$}���k
��:�戯�����5���抮��w��A|�30M	ss��W>�\l�2FjO�V�I8�΍]j��MZ��$�B��������h�˂��w��Q�7ѯ������5(�\I@B��cCv�L��>AQy��͆�*�+��X���BP�Č�����U�l��h.��(��*�p�"�C:^�һ���;~ߒ�$�v�E )���(Fxf��ߪ �]�0�L�zg���lV*�b'xYZ`���3(�z#�ƈ��T^��5M1�7f�O��r)A�SBC�<!r���Q���+���Ȗ*�@]=U���(���A��+MŃ�$W�����S3m�����[-�3�<$ez_�C��������hk���Ҵ�炬'��ET���v'�yg��$�"flz7-��w��j�4Lx�A��%��q��$�9�GE��p�ǛaZh���T!KA�J_Њ�Z�;}���H(�|9I�E��G�n+l�~	"~�gI2ΨYH;RJd��Ȥ����xw���?
�����
^��ѻ1�T�fxGw���v1�c'�^V��LGoS =�:�~�[��m.>�yE��pr��@s�#\���_G��D�:�gH������4��#����w/�F�u��d6�}�Ιt]e1�&�}��!4! β*���gB盾9-<��&����~�{�9��;���D���b�� ���r�i��RH�-�����<��h��h��ɶ&������^� ��|z���cl3lٝ�����R��]K�~�E6�f8�p�F��\��<H�y���g��{�:5Y#��gI��2�
M�!棋��N�r$k��e�5�=���7hd�O�)�j����F�NC�7O�V]AF�g��U��w�Ư�<(�W�kK2j�%���^�GӡWƵ���ݻ�(g�������<�#�v���
s6�ffb&��zT�Gy���|D�6�(cJm�ihjd��"6 9���g�p��O���<�&h]�`ڀ��۔_F�*N'��E�x�o­��i�낼�p��KxSx�°C-�V�Nj;��z�4S�����wl�`L���%܎#O��u��S��෿��W�s��L;�X'2P*�*����#�as������E��.i��\���b6�|N:�Κn{J������]%f�0�ԡ����6��f��*3�"ұ�T58+HF�?�m��ݰ:�����&��E�ᴰ�6�����{gB�Y� !x������G~��.�}^�Yx��<��}OI�����uNO&L��x�R�D0.��2;X��۱�C���S����^!�\�7OU�Ҝ\�ٕ2q�K�7O��\��e��ޑ�M��k�-D71��ngu��h:W��G��_��7\�w��,��F ��3�O�ml"?��WG{K���a�(�p�؋�dj2G��3�Q�6ߠ҈��,`�5qc�y�����.j��j�.�BZ�#�`�T�-u�GhX�i,q�=쿗.��Ue������[�l'HU�
��80<�ê�ED���r��p�c�&���7ʹ�d�̭z��¹R��1rd��c\!U����<�e�����^���}��q�;��I�1��U2I���G�.1�ԝ&����2�+�
ДP�K�]�i���=)_`W>o�0��/���\w|5�]�Q��Hjv\1IN"�q�ku�<5-���vs�Jk��z ?v@��]}�?��U	��p灌��B1��ԭ��Ֆ�m��8��ee��z\'���W��G�d�cP�;}�\�Ke�q��B7���8����������}���^���<8��J��/�/nM*�Fw"��M�T9"^!	�{�MX�n�[Tw�~�5L�.$)���a��m���f)rM�ǮkAˆv�>	�@���V��Q��"£��#���7���_,
�}��cҩ�
R���@W��Dޏl(i|�(�]���|t+��������U/o��B�	2Ԩ��5Y�b=H�$M��]w��Q�٘fV*��Q�Z"g_���{$Dj����z4�Z���
�����{���#E�C������{�2�9�O���0�M\��8�9��w�����V�/��a)���w���K�� ���ۆ�����z��,����ՁL�ե��D����z:��q��'�
:�N�k�f������q�nLY�@�pt���(��O�Y��&^|%�0z)��'*mB��[)��d���V��\��J��ԚEr�"��.Rڹ�K��g#�	��o��~P�41��vC ��)���M ��&1?o�"��F\�d��F�o�,�x�n*d��{���A������kn�2�S�BY�|�*W���|`�6ۚA\T�� j&ٻ�mNg����}4��55.�Pb}k+o�w��C�ӄF�F-yc��y2a�4Qi�	G��|J� G�P�У㤶l��ke�ҹ����cD\̎ Q�]f�1�̱��_a��O�s��� �$12䰝f������p� {��l�~v朽O�oH��=��V�E�B>�f}�A�t�E��~����A�A�Ѧ.��A�t���9�o�Z���^qޅ��|+��\%{r����׻���W����X5nW Ǯ�ֆ��@pn�~1U�(j��>��>j�;u���,әܳ�Y��I�Sز�+%iW�o�|�tec�әfr�&�c�J����b��/��.9�w��?'����YSV��Y=7�^b۶dx�+�@|���G�4o���zcyjss�($2���Hs�QVV0xd�U	>�J��\E�$`�(�����9y?��h�C5{i��e�B��(C��C,A�]�.��� �ă`s�Ԣ�8+;g3�J�m1,ȍ?�-���~��q�uW'-hmn�"�򘈒�d��>⯦I���i҃��wq���v���,;/3����=�%��V+�|ݽ~0�,���\
K@�j����"_(�0�b8�Ҁz%t�[�խ���W��;�쪇Z�v��V���"�9��n�օ���$���y`�r��n����
�pۚ��0rz��+���K�;����'��W��J��΢P�U�0�gl�XЧη��A��)�XҰ�}��Eiƈ����$8h�F�@�D"s~���ꢿX���]Pҙ7��[���)]��N���%�S�ξ]{E�)�"�xsUH{]���Xʰ����SX�N��O�U�ztA�JJ�Ug�����T�l�{Wh��5yt.>k�$E:J��$f[d�:�qE�9�Xit��坦��Qx��=���e^�[�5,גe���Wc�_�V�fD#K�}	���"4��?�Q[(�R�@���aI�h�Y(A�a��!!!�:�%4�.���VJgHy�4�7j�ݷ��H��t^FF4{qK\OR_�`�c��P�e���Za����¤����h� ����o*c�L�))��<e���l$��%v=�WU� ��q��)�K��!|�""6�dk�^��>�e=$yҡ�0�21�7V�c��"�hl�����%�GR�		��yۑ��o��uu��oX{�����Z����A�A�W����̢�c��M}g�/��L^�a�����j��u&?^c����;��d�$��@\ҽ�|@�>~>��w�Z�uL鈡�cYg��Z���"�踖+ޫ�A��n�6)�G7�\ ����X��}�6�>">���xh.&�i���s(7�\3����Ta�,��1P�����q�  8���j���]�z�66�K�ߧ�$$�V�`!Y� $��H�v��J�-��;��_��G͵Ư}LU8���n^+��P�?��|��2UkB;8��[��'�!_lz`��b����.���,h�O3P����b�1�)��
*�L��N7=�T_מקN·ʰX͇��Q�:�|�_y=���^il"^��wt���
+D'�7td��x�?����G |=�rԏ��^��VA�e��U'H���O%+�@��	P�Z6.��.�}G�}f��Tx�S;6M,w�~����탆�*�� े�~�K �K�����4�%�*H��>|�]���~���˰d`V��R����7� �'Š�M	�q3;�o��+�p㿻���m����jYY;Q>J;�z.�1����3NE_j��@P����-{k@O��Q^w�<�������$t�5�L��ɡ�v��2g �����6�=�/=�"�PIn���q�.���|��4<�X[{5E�	�֔�� U�x�=�C^�t�Į���\�M�Jp7!b�~���SN�"jT	�b��r$���bvr$��ῠ�N���-|��&�Z�N�f�h�r`����D� �h��$�zY��(��h#��$|�a��JM<�j_^�pݠ����W���
��~=́M]L�J'RBP6�1��-��W�O*aj��2���_���<�A�h]A&ϟ.�S\������*r�ɲ����/�|�ՠUV	���Y���W!��'?(�]΀!$�X��ڷgU�Y�������|�M�P���f��%�8�����$�nʜ��zQ�S+Oa�/Ö��M{����s%p�#��p>���\|2.za��Sig���S)B���� ,���5�0�fֵl����rL^`.��W���m2��BOm8T`�
���?/�\��4�>m.��A4�+L5O�82I�Υ�x�eݱt��o�<8�n�>g��c;?���o�p>����֟���.���WR<��ϧ0���L�f���
��B�}��`j�s�ǟ��(�I��+#����5�j�["��g���th�͎ �˂�{��MD�Y�2�]õԡZ?`T>��,#ۤM��B�[�a[�w�x|5��}r�N�6���/��jRE�=��Wu��S�s��*\�m��W��i'	����@ J����﹬�-�]0�ƭ�00�))�4TC�(>$:ܫ�U�d��Y�m&R0LЭ�9!ǽW5�T����+;�/i�yh�\ [��l�g�2�9&ǻ�.�� Zt��X��I�vXwD�o]��z����Σ�*�5Sy�N� ��C:RP�3��M-V�����|��Q�)v�{����3W�Q�jה�Ĵq�H�g���u�����WtJ޿O	_G�f:���?�����C��,��@�#�Z���:�n������W�V,�L<Ǘ��$��e9��xЦÈ������ֶ ���Jd��s*�$���S x`���S�Q�mI/�PphZ3"�ݥ
�H��=�l��%��-���iN�ׄܢ���ϻ�X�g@�ީ�5ŃB� �k̒�R}ǧ��>��{��UPRz�@x�a��ڈ�?�l�^����f�J�o1���+�s�Ff�������K��i����"{s�kl�UT���V�ӳ���<v����|f�54�-�"���ٱ��?�u��#	��m����i��� 1Ud��T���b{H��G\�;�L��f���6�k�W����B:��ҿ'�<9����n���/J�<p������L�����w6Ӻ�\��"��dQ*1�+N�xP�[	/~z�U9���M,]��	L2/��*��p҄�@�Q~��g��6 ����T�Bm�n�Ӡ;�M,��G�#xٜL���B����d����t�'�x@�]�F4i'\G�m%�r�A�j��hz8�%�0P�/�n\��)�l����o��0FV����/����"��T���������iF�����q�?x�m�6a	?R�_�~�R|SiU��mE(Z
�� ����-j*8����.t��2٠.aE����u�Lx�3�����zܾ���<���l#�|E���b��p�����@2t�L>o\�"Ed���tf�/F�?17����|Z�5�1^�yv��+��JygJ�x�[,&B!A� �`@��o
h#����>���=�����C�=�|����π�g��NI�C�����s�H�n^a�bY4WDP.�
Gf�æJ��A�v7{��7y��aF�]�*�.y������ٞ���M{�>��<sy�)���!y�����Q=� ����6��{Ļt�#F �J]}���:�_K��<�[�C�U	G��)�K�:�8nɑW�� ���2�iJ\_t��"H��>�%��L�_��qQF e�|�	�@����c@7{�y���9��7�͛���i�33^J?��,��F�����XMx�����ڐT��$�em���l�m]��d���t)��m7���5�C�c�NI�b��,/iĠ~���@��F�:��Q[%�U
(���m�y�j�a�^��%�4���^�E)�V�Q�����MDF����^b�+���WN���6[ȏ���N��*�ųˑb95�Y0ߠ�v~��hE�����S�]���~��q#��5Oq�s�z��'���'z��AVcT�#2�N���oE{#�����'��D"�X�D��W�@)+�ЀJ��:p��mA��Q�-��Y�&��j���E�h��W�qdh
��e�e��/~Tlٰ��$S��㿬'�Z���.��y{n,��B5Zz�vkQ�(���iy�řD���:KB�`�������'Ҏ���*���L��Q��΀��!U@:Zm�׮�p���"�pQhP9��Z�� f��n̖>`G�b/���Nd'�(�Vo�]��Bǀ�����@t�7}��n��&u-�Tq���������+���L���X���-]�؝Xw���ڥ:�/�ϕ�+ĵQ0��r>��#4�W�W����lד�*s�C
�:\m)+b2�!RC�s������*�815g�G��Y]
�O|��m��ן{�e�6ET�{
�J0f���7P�B��qYa��&��,C`c6��>��/I��}�N��:������������)�O�-�Դ��3����q���
 CYq�!n7�[�(����yc�~��-V�g���#R�ȧ$��	�u�nJ��^�G_�(L��b�}��g��k�tV�C�ׅI{]ɸ}�0�mhհ\�X�z�*�{�\��U{�҄�(�m/u]�Y��|"����]*��1�(_g;�̅���z�	�'��Ǳ]�^���@�w{]w3T��*;O����'��0.�o��T�1��L��P�����	�*IDJ+x`��ܠ NPl������	X��C���¹N��2�S��C�Lk��s����"�C4�u��T������'��Z�h'�t���{���+���O�����
��O�:�����$�G*2XXe75����i_�v	b��sD�J�[JK��?��q��E�]��N��~_M�}��S�t�ʴh�$�ՙy�)�������|Ğ� %�-�R�n*g�����@A�ɢm3^�㶄&&A���%��5y�wR�f��Uv�q�bvu3����}*���d
u�hK�����J�lu��Ѳ�
tV]���=��5+�=z���ߧ�[���B�V���q�GUi���)���ܑR;.�:Q���C�@vxI���Buɣ��j��RϾ�]�pQ��b�{�R�q<�+�-�W��¡��3����%�D�Q����-�I%�qQ��i�B`�����O_�v�15����<�8;��:$�e}n��l/x?�+/�u����AtlC�I5�B%_d�.���޽�/��<��A�F#���D|2�I_k�C�l�n���K�O*�{U��h"�i�|���`�n�����k���V��0�
����e����^�V<�����V'�`�s�t˞ׯe�b*r�d���}{����F�D��d��D@Q��ڊ"VO�b�|�գp�V�Q�W��[���`���{�8wM�6���J6D7��2�'3�6S�(�B������%�{~��Sg��=Y����%ê;i��m{/�0m� wu�W+O�k3��)�X|�o��x��H��<��i���4+�Mg���R�۰�6OiߘH]yT�t.U��~m7F�n�D��h9�0�W�.�[p)f�;ua�8�(�Xr#Fʜ��ٙo�xlQ����to�s� �{'�[�p��kN�S�/*3Oe8�2!��߱1���`�]��;���؋�����^O.qr*d�������=k��YXK��,�U��#%�5=3�DfO��C��Y������8������V��T��7���y�&��<����DV�il��lW�&���T�O�:��4�v����X�l/x���Q��JPY�#Y��=kW�}�a?s�D�`e'�6-!�8����=-hSS�/�z��P����h�݅)�����6�]�ʟd��)WU��4�6��V�^�=�I���񅠱�d�;x��%.z��`���[�m,!x���2��㌶��$>x���1��t�h]KkUυ$�F�P��	C��)�+V*0����KQ�ť�T�t�ok5?���!�_d��9B7�@��4�F��yR0�D��*�`�E&GQU���4)@T��.�^�	�lŋ�����
��s���%6�1�9(�������6q�����uˊ*Yi��\��f��6~ja���i�C�u]7�Ȼ# �XV)�lp��ޤSwV�EI�>��+���e��ow��a@E� $C�z1n��#��*o�,��`e�c	�)�ڷ��Jt����zy��N8���JϷ dfI�K�Z�O��X��bx������}����P+��l�].����9/̀�|9���D;�R�_�RN���|��Cl�����4y��E�k9q������R�Ľ���3k�6d)l/�,��&�@�Ǉ��^�ʨ��x%�7�c���'S��$���e}��ؘ�]]�O�M��U�v7bAM:	n�)���AB������=F!�B׋y�P�ÀW��"o��Y��+����A
T�"����hQ�X��'�Ǐ*Ť�ݰ��u��[<5� �I
�}�dŸţjRR]��"����l;Y+k�
W����2�G����o����\������{Ç�87���e
�!b�д=��B�C�i����2���9u��,֖�	�tIҋ�̞���p+m�-f4�^��a���q�*�c!)׮����G�!�,hZ��i���U�jS!���N)}U���2���@��=�.�4�kl�>N�c
M�k��NVQ��c����TYW�p�͐�s�	�d7b����O^���(ŝRg/H0��a�6���`���!4.�O���@`�#�t��QW��s��?\s*����FoȰR�암�����3�t��}_g(g��
�K��:�O�� R˕�8t��9z�#S
�.?$�����S��5BA7.K�����}h\c�E������ɵe&!�������츎	�G@R���$��2��p���L��Y�U.F4n����l�R���,��Og#�>4�gr�b���XJ���*㞖̂:JM�}J��IE��}��Y���]��%w���&W"���N�xir][�V�+���ʴ�׋#{M����oS?�:���L����I�ÿ^��O���o���9�����~����7��ZZA��-��62�4k5�#��@�W9s�Y����Fo$�&�E�1����:aT��KЋ<u��}��ó*A1ijާ��X��i�o��uP��3��c���"o��*¹;溜k1���� O�ƃvDR���>}�����:O:#3����fJ#�%ۅbm���G�`�ksD���G��ሤ�-����!,���,����NN��XǦ"���/������
ē���:�~�䜏ɽ)~~���0�5[U���wx���ϲ�6T�`�k{��a�R^��҇:'��T������
+����3/d�e��3�qQ���j�۲}��b��z�8v�!;#4�<h俌}�y,_�Σ���Vgr�ݧ%)�;C�����H��GP��2�T[Z����[���%��EJ��魫�e�Ŝ�m�Kx���!�g�k*j�X1��7?��� ]+-t��r��%�rc�":���(u���|r�{&T��v�y�x
7Ԅ�
e���4��y��3��−��:�nm��ۡ}a3�	-ԕ�)��bS8�����j�z=�H�������Ev�����O�;p�f��R}�0�����L�&��xa6j�����&����G'A"R������I��
�wHׇj�w�C�%��W>���##���ܦ�<t�I<"�!XF)&m� �GSnpU#܍>ا�_-��j� �n_~�Y�Y���1��w��}9��Y��tP��kYJ���� 7��1�U���$}�H_<U-���Ƣϒ5�.��77A���Н=Rg�i�2�*��1t�,�^����q�r�6���*k��l@�Ῐ�ސƗ�i!�ig�x��	b�ʈ�w���M�bE�=�Y4�.�1�Ղ�5��F���@>��ہv���x�`*�T�MGRIH�HC���YM!3�2�����S[1�D�� ��@{�@o2�GI T
"���?1�R�z�QY�.��Y.2B��2(p�+?,Ҁ�0�=�
�	�&%M�-#�#lр ��C^O�wz�ÃRi�����T>��,��o�g�x߰�-�	�{�	ܮ	f���6gY�})Q�������On�������'J����)��|bܩ��5`Cp��+Ē9��Z����z`r����������1<��Q��Y��$ �+���Ϫ(6�u߯��KW��}�iǜ:/$(�j~�@��P�8�$ ^���Lh���¿c��H�6���:����oe`���#�P�<Si3v�ie�~�=���3�c��%�X$������IS�3�Q��W��if�_��O�6����K'㼴���L��MV5=E���n���ѱ�S��3tx&uD:
ĸ5�ޙ6XOo�C���i�V| H.�F��A=����!%jq��U�4��R��E��GR{�cS�G'W��1Ą�hJ�)4��$8�p"� �B����C	���t`͊K,�
��Q^���$�������&�،�`T�e~�J3ǈs��@�!y[��y:�����VE�`w����A�E�d�E4fw��g�숂�v�l-��~��J%$;Zx6�O#��V�I%�����ϳ��A��$���?�.�o�F>��O"���Rio=b�+�L��b�~& �Q�y�]������ۭO�����=K�	�W��S�]$�2��Z>�C��It���&&�C��^�4͜Ӎ�h��%Pws{@�<OL������d�6���y;蘮�^����t,lu%$<~/xb7X&*��5T�������r6ݫ�75�6¹	��J�蜌F^:ﻻ�q���ш�n��]����pFHG��ex���q��d���'�Z+c��듳f$A+9ޘ�\GE�"��j�TY�B��;lJ!���8	�Jw����j���T��{"�@��S^�V%�Y%��FaB?���~ T|�"R��l{:,�R��K�Ɛ���jAlV��*ze�@�*�q�ϐ�5�d�"��l�HN�zg�1TU\��J=K6d)T�/v�R&�6����!W;��:Rb�އ�HGc��?�~��_�LΝq��o�z�5��^��C=�����j�w:�E�]��%t����=-�����������K�l��#���f�D2,F����n7i�W1s�R��>�Z�.[�^Cf��'�[�C����u1��Ox����Ӥ�����v�����<-CZ�s:6)�y�sZ�(`BbQs�8M�<"�[��D����ܦ�q7��m�B�+�l��E�;����D�	߿JG���n�>6��vd��s��i�'mg{x��b0)|�ٹ� 98�������ތ�,j�W���֭o�`��(m#r������(��2�!�C�q�i���]l�*���,�
�j�)O=�F�Ǒ�|�F<~u_�Y����e�<���X�R�jZ�
�8����-)��i-����K/��~fb3D���]��k/#����A����&��r�ca@C��w�~J�����-;P��sxE7�hˑG"�u1���y�QO�^e�ڇ[�1�C�Ewl_�J7)/����IL��5<�>��(���9I����D�r��|�w�k|6\�ҽ����*�M���:P*����x�愂J�a̦�����]����O�o��5ͺ�ų�)��������Q(���"���c�BR��$y7�:J?>��?>��`���J���.`Y�a�	�K�	#�ˊ�%׳��o � ��F�(a�PM��\V�N|�ot
�`�Zp��e�c�4>9+/ :��'�C���Y��r�&	�k}�����4�~���RP�+���W �˔B�I^�gT朿<�gֈ_��D�(����4T��cn��K�d������U��|B�\�|G���T-q����gb���x�.N�@�Z֐�*���z{�_��7���
��!�.Ek����)�+؞/#w�~�~o_��߻���ރ$��۫��:jF�ڋ��F9��3c
��E�/I4�Tm�z���]I8�V���泻S��忶�{�E̓�9�M�V�U�r8B�4��V9A>�4b%fK��Z�h��ĉ&<�9�Y������T�4��C�j
��r�8���q��	�f
����D����Q{d@r�t��4��k��O8��w�4�W��3^�]�+�wUX]��2��1R��l2o̻H�}^�<�1͗�iĕ�Q���c����G4�QS�ͧ���c
��L�.�R,(�Լ����x�\�jV�Uy�V\�ր��ȣؒy��i�O+B�D���.��JYA��^��`�}�}7����¥)gy��8:���ݜ���A1�ApU딦��F����%Ǫ��/��6���.��p�z
õ��a��>��0�N��z������^�V�֚��GN4k�{���!�v(���H��i{��lQ��c�9v�Y���H��B�s�Xq�yc�3J�7ы��� �K����,P�J����0�E��I��D��~ץ;*;���2��5�B'�l��|>Q�1!]Nw�h��0SR��6�B�#�>���ϛ�YQ-��	��%,w!��k�:	YGPXR.�CR^���`.!eԕ�"P��3�C��	��_ENVQ��=U%(��p/�Ĥk�"W]��	SX�6W�<)\G>fg�5�� �%��}C�ΰ��)�5V)T��'GJ$@$R������!���Ƒm�O�%vH�T�`_d��}F�N��/Zq�d�Ǖ�S��D|�*�+y�b�@���<,����P[y���W��E
�P�i8�!Z0����
儖5�8b'���]�i����JQ���VO��y���^�\�]1u��W���g;yd�K��'#��D\t��P��P�Zfi7]@�cܡXb��K��x�F�#^��@=1��RX�+~��:�e9ݟ�"����طDeM�TSg�U��5d��W�J�9�^T	z��_��8�TcA`�3̇v�|��y�"�ߚ/8eJ����(,���c�������oA}�k1
LL�嚦�'�N���7�UTliIVI�PL��1��@�
�V��	g�ȽC���*��w=�V]B7�
T��GCJ�r^��º�(2_j�?q)z��B�=0Ϛ/j��p�4�+�Ha<z���a(4(�PYs\�r��$?ս��T�XE1*�͖@}�Bk��5�HD���� j�mV���:yl�P��]M[�)H6lԠ缙��:i�A�6�yp|�B&B�����qă^e��L7��v���7�@@7�B�b�ohqN&;�W�F��9��(�Pٴ��C�힅:��st�]u��al���oF9�y����}Q+Z~YIUiJe�E��k��"�Z�5�
�U��f�,wxP_�I"k�{�qI0䵸�����ew�]���uh�R����6�#_X�J�Wg�00��H������=PL��2�]�)Q�'DcAAح�J��GI󅮖���� 흒@R�t_�R��?�y�fK���i6ù� �}�58��V��`ͷ�����w�:(끢#)\�+�B��!$��	H� {-�$���+�܀P<�iR���5U��iKv�c.lYVt���_ӣ8v�>+��|���U�O��r�����������dg9j1Je�O^[!�|Z�sD���8Ρ�g���-l�`#��Y�8��X�`�q�܋: ؚ�9+F����ns4����]BM�a1^S�CO*W��-�"��D&?j��^ݰ���C�b/��A�y��: �1J�{�9�CH���V�����i3*�"ih��Lo����ww���gzJ]�c=紉��Ӄ�i�i�+����!����c�� ��1�w���%E��ڠs2�B�66���o.x��&͍;�d4�-� �(���2������ͱX�� 8@�HCU��(2[�[q&�,^�s���ha	����jf��b�R��It�� �t<�7�(�a_�2*�����S@�Q�m�/-{�*$M����¬Q\��g&����wյ8v��'N����g����`
���w%^�E��H�=����t�����MCM/X���JY/��i�sL_��n�.l��P-d}��c'���îV��h9�W�����C.C�HT'�GR~QNM�p��{���>��w�!���;H��W��;�C�Ǵ��C=��T��Ч���/�.���Ғ5	:�ސ@L�u�3a(
@c���1�
?��@��16���+���,K�m
fad^+��o��D΃�4R"��Č�����bN�6ƴ��܍�),' �7����+�e�� �Wd�ԛ)p[B���*�~���Az=^�uI"�(�j`�%g�輩Ew�݀Ѣ��"B�MQ =���=+zU��3<��3d�G���3Ij:	g򫯙AF'V�;Gw]PJZ%�;�57���:)C*��OH�`p���M��u	���EQ�:�S��T ��S�������N�8��q�g8���

f�x�ڋ��ol��LVL��������T�v��|���K�D�}�띁�t�����i��.B���gu�ﲣ:i�m���r7��z�8!^�7���ඁ�,���\��;H������e�2��^��+lg�0lM���!$���v�ҿX�5u�I��l&��i���i���l�/F�ZH��D�����6��!bJԑ�m�; z�c:��S�U��nhp��[q�+�^3X�� A��n�n�|XT{�9每��SN٤0�w�Dr�f�7rY��l�6Q,�[�Z�.G#<�����S)�X]\�yB�I�kfp�� P��3�(C�f(�D6[kU�j�A�_�Ȓx�Lo{^�F�����[��"�|!��Ѳ7�s�R{��l��t���t,�"0�Z�EIt7�qY�� �0�dx9�Ca�8�s�˯���:��Ǟl�~f�3��*sg@�Cm�
ˤ��R<쩰���y\���+w�'�F����M�˳����W	Y��⨿0���w����_�NH��r�ܑ�1S!X\t��}�DГ���{��x��Ճs�e��/fnNq���H]t'D)x���[b-�����]p��P*���Q+ar?s�͟���1����F��	�< �Yؽ<���c�����@v�~�y::��J>(Z�8O����5N;���		|3}�
��S�I
��"�/E��+���B�鴰��J+�۲�m�����7h�JH���<�[���]�Zmu*/��A�_p�K�r��	1�?�L�T��fnG�]�?S�cES�MCaҺ��z��ΕXF�����n�ĳ�!]�#���5�3��U��ך�Y+*�)'�7Ĭ��<	4������CO��2�
�σxØssQ��|���8Y&C�H����[� �I�@4�z�vޟY�r���N�0�n��p�F�J���Dx]�eT]�l��S�_�Z�"�w����=.��Y>p\oIZ��:m I;�ȱ3���.������XGf��SM˰�D�s�m}E:E������j�ņ��љ��s���Y��&�-3
]�]�<���G�9�x��vD���J�� .�H��@낥�i" V�|t����F��g��E6�HԷ���D��G�|6���Ww?�a$]0�"S,���X\�i?�W�\�9aDK���1ok;�{qsg�������J��%AA�����Kj6��USė�Qo�������������|����A+���%$(��u�ݿ��q<h�D�����P�������zC+i�D�u��l7A� 
%��ލ`rNr<\���rҐ_G�P\H�9_h��Ih<���%��6f�Q@��-y`�OyUc�;��S��x����P3��h����Ȱ�.U��h���Ɉ��$_�
��@^!�+�qB�܅Y<�ҁ�*)�õ��l����X�d���qT����+��}�u���H��IT��p�h�����GA�9������X��/pB1�޸bM~<mmܴ����D��ܒ	){�p�F���z��;��.�l���`��H@#gF};C��i���w�WL���k��u�:�x*����0�e�e+$��#��c��Y�=֧��ԧ�Cv����u�������R�8�!3�v�V:��'�2 6C��լ٧g�C��Je�������YV�Z��}�%�K�E���Mct��.9Ug����t���tp%�$����$63��*y����/�R��+4"!�O�)]$�Dfxiq�mT9��/eg5�5��:yO�so}D�=*$�[����n:��pJ��gUW�(9�&�����Zue�q����}}X�Ǝc�:nv>s��H܈b`�2B�Qq��{�*��P �[ �����8�6?��(r�厾����p��B��}`�� u�Y{�j�:i.�;���>s��?D����{6�H�R�S�F�Ϸ	)ۂeLsF�0\GB^`�)��O%��No"
���.�R���V$I)��=F���W������&М;^o��0A����X��^��,�!�g���0���=�-D��``��]�Y>W�9L��[t�.����Hq���i���[�r}v����Se�-��7�}-	��*��s�H��	n�g�8�ġ%�@/L�G_�����Uo۫��X��V�IG����YVv�ߒ�Z^�e�7O%�|8K���I�\�F*�S�3(sd��<OhM�
I���x���_ �1v��0ԋuAh����-v̅�`��G�q��xF��j^S�А��Iw ,[@�a�\����:<���@�j:3)�����?y��1��OB!�&x�q���f����-�V᭣6y�W��%�����(~ rk yَ1���Ch.鹦�=qJ5�<{�^#o�:U���C��1N���%B���7�b<�C�j��{ �v��T�F�6�P%+�a�5�󉽔3�S��F��xC� �..�#5�vd�*<��V�
�>��'a���%9�`Z���4p���Q�N�@l��v����+�*�Ȩ�u�DU����ԙ�G��p	R�"����� ���<A�f�ƛ�H$�@hV�ݡ��O"�r�����4���dcy;&*a����t�⟃���W���Q_�u �� ������jż��0� T��X΄붥��#hB�_��p�d��CΘ&J�!AY�#>8s�:������9,Z�o�g�����%���T����> �;�%����Џ*%��/M�,uxo�2ё�d�e�ٰՅܬT�^ڠ4�s��;����~_��
_��08��
��:��ќ��%�8�y�g����b��
rڂ�G�l�R��ȯ�����"a}Ѐ��noN$45K�KY�x|�\ք"<�du�Y�79EmSd=������{K��qoSses��Ѹ�JȆ��b�%�K�42��o)8�m#����K(2������3�~�Z-l��b��L�X�t{�R}��C��~�.�s�$�W�J�^�v�R �������_ᙱ4�))�(�]1K2wm˫9a�z~��#6a ���ʳ����KJ"D���n���\��F�8q�[I��MH��T/����ʢ`������!}B��n`Xix�I�5Y�c:/�X���])��9�9F�K�ߚF)���5�"Naq�fS"_0Q��l4�(Z=x���K5�z���y�F��k��U ���o��el�q9�EP��:f�WOtK4�6��{�WhO)#�m�C��������Yi?���>t9|��o\���&C�蒗龣W�4`)�3�Cr'���%rT���?yɌe�W,ƓxrH�毘�BχP	tҩ�}����cQo���/��Vψ2<�3S,.rN��ܴ
u�i�����r&��y��d;�̡H�-oe,ﱑ|��v�F�ԯ���R�3�ҸD�;�n�J�b�� j�ʉ�gl���t�Vj#�4�$=����2��	<@�X$�y �X��"�_���wB㾰K��4�2U�VdZ�U'L��~�ł���#'��~��J���K6��PA��zLD�������:H�R�8����f���4�s�`Q!�<@AC`� ������>f���JYg�6�Yt�w��Z���I��μ��
u4��W��	y���
\��7`=��,X;*%�Ýd�O$	zKáP�����m���G�BA���(	gb>�%�ٳn� z�����vE-9�t��fc`cn�`Ȥh��C����T��H���[�3��/1����􃹬�K��s��ޏ,g`[�����\���^�;������S��㥱0R�C�,C��u����r�%	�o$�H=��{ey�6�h|����6��:�aڅ5^؞+��.A| �O���Ŭ T�WJ�F���4�+�K�!�8����`|�����\O�^X����@t/Og��ɬ����E%&A~��rm�����e�DV(b �栚�\Q,S��u�Kk��[	^���ċ!%t��6��/�k�C�.�IM�=66��x2�>:5.a�A����sB^��S�������l;�����	�X�t۴�v�3` �8�T}���W������2�z����ۼ���33P�7����f�vb�/��r�|�d'<m�NLS����Tx�ځe���W��M����4�h���Y�+�a�4K~��z�+M���K�'|�
�X�ӣ��E������ԇ�N�7d����t��R�5)p�V8�&)��ȧ�(R�EW�z���^Mde��e�
�˵��u�tG�V��B�/k4���߆�~������lj�p?R�[���猸���N���N�H�����8��n�M����m�/}b-�bZ,�k�B!
��ko`!�:s��}]�+Y|R���R��L�y�0L�N-�5[�{z�JU���2����,	�BtP�*G�#g,�h��1�o��GS���1?;�;�-3]ߡ�I%RF3�8C�٭�F^��Eg�lx�}Dc���#n�7{�Gɝ�u��*E#�"f���,M�
F^|�-����f�֦�Y��*��~���)b�rMK���nіE4�q�/�D�'*�#�I�Ǧ�3�G�ư�������H.���|�{��R�.���H���?��]D�zd��n�E�T�	{�\ɤ�K"u��Sc:�fL�eÝ̻�qD��o^�M��p��k�0\{�����p1KM��51��;����t!'}�N�䎬�F���#Ϛ���	����7�$D��Í?l*Ѩ&��u�\ׄ!�!�N����+)����UfH6j��żmc�޽���[^Z�L�+�-��=��A����6(�M(����攮�E&u��~��}1��B*1K��Kw�ZT���1�:a�pLBZ٘O�w�w��Sx��{�3�xq=�ʹ(�H�)��\c���o���#��h�M�AM�G ��G�$$Z1���*�G��v��y6���%LEuΫ/�_�
d�He)R��f�?�wO:Q��La�@BX��Q��SF 民/���d��5kj���o3�V�ǧ?����ר<�B���A����5���n9�!�^��F�[i7G#�QwH���H��H�j���V�J��ĺD"��V�0��4��5����z�[�+F~����T홁�l^Ʊ�����L�؉����,����iU<�Q�a��zn��lC��/bL���+�!�p-$�ً\����!_�"}�j�ðZ��R�E_�`�+����<)�$u��؂�X��i6O���Jl)�:p�pe+�.F!X�`\ʦ�8a�˳)��1"ѝ�W'Y�bpݨ�jh)49l�����KevB�j�)f]y�p����N�������8���8�0�U�dք��F�^��j�����a�QO�e��wnt�4�c<������r?D��( >2ߴ���ա�*���6�h>���l���5���V�޿���6`g;̆s��z��W�<	"��0�'Z�ϑ�e�H7���𭨌
x#��Ӵ�t�q��oo
�.F�؜J�E���w�]����������,�R���8%Q��Юೀ1BQ@��;�~���8�̐KPX �j���CBg<��;�9������g�Q�!>���V���
���K2��یӄ��㣌��xg@=�W���b��)a��B� 4�C�Z���鶈Ľ�N���������]<���"
)6�>@�}s�{�r%R���+�B�AW
��Q����|�.�l7�o�DcP����[�tr�m���9�6�d᧸�2f�:�<|�^��jT�i#��e.��k��A��,���M�������v��DM�z��NI	�I3ٱd�q��m]��Ӝ۳ YP�,�Tv���!�4IIE�z� �`�M�b��?*h�``kӐ�=�;(�9y��fȝ��>Ä�.-%��������C3�)�̤��fM�Y ez>�]�Fw\X_yFUڪ���	2�	1�nY���V����q=�HB]�+M�L*m����K����ie��zч��ˤ�h#�{�uD�(SL���)ۘ��J�=ď? S5����V�g�I��{�`�Y�NY���R�B�/��|���hP�0x��v��y�Bo��S�v���}3[\�"�4B/�[{e⑛�j��^���ސ#*K'�v�ZGx�A�)�y�7��\�J��xZ�k���*�h�͹��aj�@����H�P3><�yH?���N��5<��ە'��?�����9���sg�(�eG�b�r�\:�,. �����=ٝ���ه0a�Y�Z=�b��6�*�n�4݉UX�Ax\/U�0���N���%��-M�'�n_��ltäڽ[N3��e��t_҃�~�Je}Q�jzP7���F�?(��L��MT���j7��s���8��eƍ�_�H&�_]}@}5�q���lWX�Z�-ؖ�_��[`�T���!t����e�EN#Vo�?�<��y���ױ~�RA�����e�w���zq�=��¬�WY��{��P���1\��E����af�	>�=��!��M}
�yY
�B���?�KDgG�pCG�w}�I�LR��Mwа&I���n��տ�Wv�t�3᫖���ҙx\�����&����]�Xd^s�b������-[��=�&0�E�F|ҩd@�����G��F�����#R�uE�:�'��酽��'A��(�Ca�Ț�72��!��� �� %���L\t��E⑼ �쪬|ң��f�j��4C�yD*�EB㨣��/3R�_]�l��r:W�����.�Qh�5�x��E�2KA"A>B��"�|�b�}�ɡ��;Bդ�����.��Ձ�e؍�����A����q�3�R0���[>Ƚ83jcLF-B["kַ�G�宲�EE���=;

��fχ1�f`�r�*�֞�N�A��ʈB��漻b�t����C����W��z�/��{|B?_Z5Z�h�4��-*Ks��b >�Iw��C1�8���Y@
AA9_���r��lPٺ5~�S���������ʲ�|��uۣ,�\$u�`j���[%�^�1J�\�2�Քp3�?��ҳ���w�;�ԟ�?�ȰSK_T���t���d{Ϊ:0�i>�*��f�{�5�� q_�/|1���a;����g[�^�vh�lk�(��5�:�o5�&q�E�:-��\��|��/%���k�G?�'o�&J3Z&DG�
�t�»v��:oSIaj�&*��G��=BO�`"�#é��1��yM�;����\ �M2�	V�W���j��pe�Ҥ2�ʉ\�Hw�9����
C�2se�*� �g�u���u�[ �4�o��N鏭W�,8�7$Z`@� �̶h�"����]z#�qy���=�|��'�4���n���eL0
�u&*�����FS�6��U{\� �������Pê�2�s@��� �&�O84��Ժ�r��OfW�����đ�W�+�i��H"w�&�K_�6Uru=f��Yh��(�	cE��p�-��u���^��K��;���^�eVI�	a'��X�?MT�ƥ���¶����W�X� �=N��Y�k�m�*ܹ���Tj ���ϋ1��Й�m
��̾��/'���s����:�.�K� tא�vt�^z�U˳(tP��^l?���D1����%M�𨴇��Y��y+��k����*w͠d�t�_�ޞ|�!�y�z
��E�
\��� 1T���78T��m1&�L!��O7N���YF�^�Ð���\:�v��F�\
@K�h/%�,�íN�H�U'ɟ��g�j�"��tc�[�Q7��yj���=G`];��%ş(�|k��wX[��Cį�܂p/^F[�?.R��x)��|NXS�gN�w9]y@�bmD����"�,7X:�.�Ƒ\bT"�)��yP�������Y ���,�7�����0C'�	��SAd%�S�ק��>��Y� �6��qd����GJ�6j(�Yz�Nt���R	xf���^�r�Ҟ>����`_�l�Q;L����ϩM�)Xw�h���3��:o�u�ԓO�A	�\^l����mQv���=G�a?.�����'�j��<�����vzpVR{���W�p�SOcd��9ʟ&�h�^Ѐ���c\r_Z����+��W�ʐ:�����!\����]6�$i�o�]�>�����+���ü��؟�ޥ%ٸ�b�JU����L4�=� �S���2�S������SCk( ����O��Vk�c�}t���/�
��'���Kb ,fD��"po]_�.������bt����F�S�֪%4 y?j�<q�D�����4�����mX>�=��O����E.ge�y6��T�G9��c�Yd�<-��W�s]�5��!\c\k#ڈ�ͺ��ۨ��_�7���@�� F�\{c#�!��+�
m�v�$��O�<u��R��W���58���>|v5T�dL�� ӯF��M�녗�9��T�r_4��|y�����g�VP��2m����C��c�p��ʗ]��HH�<<��I�y5RI߱[;�n�����9��,Wd������u���+,���6=NW���w�ع?��.ًm�Uq)���%p��Re��R�%��2�%��6���z���c�����u��."��glzf��Û���fHw �O�I�v�z� {��	�}�@�Di�J�j��?1^"1>�i)/V8�~�:�*�n)�aM�ʹp����"AڛJ9�~�<T�P�����{�Ғҳk�4T��-M��i��è��lz;�W�J�����w�P]��ǁf ��4-��[�p�E��8�T��Fj1�>��.��0�3�:y9��Y�a#�r��&����/E!w���sȰTT��D QT	�ͶSg-�KKRj�P`1L�-�˂It��\���{��ztQmߘ�&8 <��$<� 
H�^�pn$じ�Zx� 5f_��i=?�iWV_�t��7�����l�ϥ�
�)��-}�3�nl��1VҪ垏�(P<u(`M���v��>]U���66�iV�s���HI1������R��.���X�u��[+�Y��Y��J��i�6�]0�wh �!=�����z�����;A>��c���'&�Y������_�IZͣ��(�[�Rk�R)�.j?���y6�R����3V�MD�?_����g�d�&Jb�g5�7c�K�I�SqU
�H��KJ�^��j���d�D��_;��djϒ��H�GUY'��������*�)���D����5.��I��rE>����Ҟp7��Op���U�/�\V��]�Q�������>�/v��t��k��btr&X�Jk��`�!g��w��e�2FN���X���]c���W��1��7�T��jޥZ,5t�,(��4���p�<kVzx#�U�m-��3	(%�;A ����w�+��K�9��P�Ԑ�c�B������xk���ܺ�'�W`��
�װa��,��L�=@���j?��s���L�]�o�P3�8u*w�c�ғ�	��f���z�e��(̙��׸T��&?5C,�HP�k*l�����|��1y�
�@ԛ	7_���U�zF\ ÕRD���<7$�8R1#)��*��8遄��M�� ;6xm$�X��
�2��߫%|�@�D�pj>�bV�4��d
��V��W������DLl�D�!�;�l��K��hZM���"���<�{�U����P��_!�eb3�#针%`Θ�ۃ��<y�.t*�栵�0Fio�i��"����x�4�<�3���O�Y~��`ޣV$a� K���?��\������`�`p����C��,{��/;�A��������;*M>j�.՘��!CSQ����sAOo�8V�j�pM�-�U��~���.3[G�������?~p�`E ���m,j���Q�Z���N͎��+��4�oʫF:������.��X$�k��F����6���_�S`t)?|)��P�ֱ��r[;�9L]^��8�e	�NT����e#$�;�Å�T�޿�t?�~���M�����
�1����|��b�.�rt8��I�a�T�uƼ�|�x}B��۔��m���"@��4 n�U���L���f��7�+�Ų�n�����i(�ִ��E�D�S�I��2~�����RV���;.�v1t�Y�J��/ߓaoK�,ݲ¯8��E�zr�{�C�N�K����2{�M ��d�E��~4���qqy�x=���uK:��[S��$�Bl�ɡEX�"�S��X�'	��Vv'Z5�����AOwd�ǰ�|t��1�f~էĳ�C]�`©�.���os��e���Q��-����ү��G>�-x���6Y[<A7.̶��}�;#T�y9A�<�l�'��XZ�V��=jt�/�xxSw[ �؉�i��2���`qק�s�A���ֵ�>"��9�ƨ�PP��/�9:�&$���N6��fw�j:"�1��XQ=;9�
�K�sl[��
��ǁ�=.fQ�܂ĉq���"�S��.�#S��	�x0h�'�̬&�a$E�m��j���Ȃ��Q����
l���A�+OY]��#؅�U��;	��q�¿�w�J�iQi��5J� -��psB���'�H'bQ��ЖB[
�Q�-#�b��ܗ��_T
�����w���P3��^>�L�yf縤#k���$bY�^_�s�R���#���/RI�}���@�'���ot�|���� ��y���\밪k[�Y'�I�/+��'���l��b{,�]��{a��ۥ2�dZ�M(�Ui�=�g��_ѻ]� �:~Px`h�����7���; � <z?�!΄��"F)�?��@J���6q��%t����
��N,����	�"�&/, �Pq�vwl<�;��,�U����c�;e\��7���+�m��b"6|���)��>�B�H_��	��|�pQ���ک�ʰӇ�����/Gq;�MqB�Q�b
���?�;Sس�|ς&<��{%W�t�i���N|��wY#��5�R�I�<�S;��慻���'ٷ]m@st ��|�d�:3kCնx�5X��B$_�d�/*o���ޞ�>�]�;�����+����� 8�&W3Ժ	. ��=y�8�J!�r�]�x�el8��9��1� >��B��j`q�R����� s�j	v��Цj�2��E)q����~h��u��eCE8j�h�hG�\E���MJ�A1i�=ޚWͧ�@��d���%�����fY��D*(�Og�X]ڔ���ذ�\�"�~�K��Yj+!,w����d�zO�	E��|������TALZ5�5 ���\Lv��Ue��EGeS�֍�m��'������R�w��~k��w՜���@�v��^jQ�7�:����B���EU_��~/�^�q�uU2�qh�A��L	 ��_(Ha�*�G;$�dZ�y��Y٧�p}-gM�|�Q��229ez>�	Cy��zA�i�j���mQ��a�Oζ���Ӂ7c����)��)'L�;��fz�I�Rmc／9���3D�W8s�,ǵ��e�U���ځ�3���7���̮7���(B��Ԡ}0�vø��_UZz,�B]����+��
��Z!~�b׀�y�&SKz�-�!�#�_��X�A��6�$�������e���;�e=��T��+"��o`p�=Jh!Ri�}֘پ���<���}�9_�V��?��$���T��%��V���Pe�%��AN�����4^G݃ ��ڱ:p6m����dn�h�-C��	J�Hx��Ў^Ƿ�e��Gdo,�|�;fw޹���Ѹ�a8T��D�Es���/1&D=�=�H����\��!Cӝ�ҳͬ�6%%��e��k�����G]A	;w�|�~���̳�k�T���C�?�Vr�등�⮓V=^��Y��+jq�o��ϔ?��H�[��%��z�4��S��aY�^	t@sB�0����ӄ��ݙS�u�����"7@-5�ҁ24�!�0���x������p~��~;�����v���F��"���$W1QVI��P�@v�Pܐc���nZ���H�ܳ�v> /�r�(#Q�{�Y��A�}�B�r��/>#M�=��(�@�Q^R��gі������DsJt�||UK�?�_0��-�|��^��t��*�V�x��O����*���g�����K @n~:���M�����Q�b��
IV�G�
�_Zu��\�
�H�p�n1��mpT�z�Ɯ۫��0����UN-�f������ñG����H�^���
�A� ��%j�ە6&�g8�0 �k��4�r��y�e��@�ů��C��<����ʱ9�ޯ�r�	�;�o��-�+{B/.6+AoK|�a7{kHa̒u��$9��)�^�<�[�K�4�Y�f����אW�UhC���Q��/��%�p�*42�c�wT��/���{ϯD#pl��hX�u�mG@��_(�C;ih���q��+ZJ% �I)�{\���D�ǱMZ F���:YqE�J�?b�dH帞��kh��o��'z������iŴ�R�N>�>�N0t�h�E܆��������ޓ�nP�7Q�����p�a٧�Y�6X�H���T���x��Xs1ɒ���i�S[|�V��pR]�g�o]ݡ��u��52���g���k�Ly�<!i6b�\��H�7QwהG�?`��\Z�C�fP��[ע��ch�໳<!|��}�}��g�`�N&��m�{/T|��F0:��ȴ�}���Y	E�9u\VB�<'��?�?9��&dA_'#S��,u�2�����_���\\�;���A|��J&rI���I��;��p��c=w��h�\\G��7S"�����mO��:�`�!}Eҝ��lݨ_�'��@�mbC��T�9^ֻ���a�T�*ߡs5�TͻIB���/�к,.��?&����3�Ȋ��|��{�Q�q<f�6Áh[���P{�����S�7q��{�&^Yb��42�@8���=F45�U(.����ٔ.�u�'��]�~*o�^��k
<��N�(M�_��y��Z�d�S�q����Uх@��}Q�`��L"�]D��cڥ����x(~�u�����[a�س{�{�Q�1�����R7t�����h�H���d2�6��pJ�Q��c ���*��U���n,�������|���D	yY-*�&N&�'�]��/��9���م[p��	J�4�s|&SP�S�����:�@w�H���(����(W'�w�؆f�j�}���:K��%?�V^2��pX�`�/0w�$/'Acק�V��Y� ��2G�=d�WT�3n'�^��L}���y5G�m��ݛe���|���<��N���7q�Twͯ��ڥ6\�T�6ֈ���_VE��Ik@^�u�j��W��M�ʏ��,Ee �d��7y��8����,#Io����v����	����V�zK�-�������N1�F�{��.���*U��NBN�db�}�JXn�F��S�2�(BY���)�/���������0RE-�}��3�,d�%[o賛Sj�޽ֽ�B�ģ��d��qK��F+VT�¯�8�����&�xc���<�m��̑b?�I�i���Nj}�Ox���}�-�Wl<��WX��0���R%l��A;O�gć�����h���Z�5},��,Df���gZ森R������,�����}���h.�P��n�����8���-���c�Up$\ Ĩ#x�m����&j_����;��||��/��~(�"ļkhc�Ԝ��Ȑ���F'�a]�lꢉO�7���J<��(�H�4Y�O0�#`����8g��@���y���7�s��(����������+X����=3�@L�����aI�� !#�/'��ř�+
�o�`�4�{�3%d�_�ݱ�}�U���K?����"he$viޭ�%���}����S@��ç�+ы��Vyz��b���[�3�R�` �7����.rMiZÔ���@Q#�_^�*�,��y��0�%��wl��p��L�f���ur��2 ���Ĩ��#��9��omK�C��[�x�n҉;��)�S�@��U(E#��8 �׀|�p�/fф��H��eF��_�����-�T����7��WFѻ�-���
�x��W���դ�T.D	���m��rR�D����� +���"j��9�+��}4���r��a�� u1^(�˴`<4Y���f�7���a:�ʁ=�J]:�p�p\-��$�Gj�9c�:S!)���>��vZ�ۙ��{����٩�3�0��?yN�YFX������dFR�u�W[�DıSkP|"���=5	�����_mb��It�d�B���+,es1JF��0[���_́
�� �-�Aw��+��+�T�ѝw�����U���G�,`���ʻ�җ�6�`�}e��n��e ��L>N�|����P��j��j��Ix���t:g�R��W��b̖���-��9� "�9Qخ��d)G��a�m�}F���R㉓SL1������N�{��ǈ��2-{�6�7I����5$�z�P�~�r�8�`o}��!���qr);�bL��-��9�B��&�������c(��A؄��D}s+?����W�e&����=����BJ�i_�uY<�ғ;
\I�vߞ�f��ɸ�W´chg����>���ne�����K7`��a�i�[�T�9V8M���M\0N��M��'���Ā�r;~-�)\�5@ً	�R�ci�}1}5��z��("0f��5�w�����<ɨ��jZ�3L\��4}p<@�����n��X��{�hr/
�c�?C����F�K�����S%����Og�ʄ�$�N^{Y�G,B��)�_o�T���o:�l,�M嵂Z\d�4v�Ke�V���]O,���z��gU>�o��L�5f��2?�\:�oߋ�x�Pf����Js�S��ǫ�lRsF��2L����_�����z����7C�E7Z��2�6���ت��	�ҏ�@����Z��f����r2��hH`�D�M��
� #�  ��F�Q�#Dj@�,;�l�4Z���G���b�ƣ��k�M���)f��<�1,�9Vp�,7i�-�����A<���'��A~6�-�a��AC� �Ͳ~�_#�_��:�O�ݼ��A�*rlK-�Cv�	�v���W���%��+4o#�2��DL?A��M�j\�u�P��~}��&8P�����d-�GlF��*4��M�A�Gt�kqX�JM��ﵼC�[1˾�v�ȊD����坒�,9��?}K��LV?5�0Ȳ3>��'һg�����L�~�$J"�x'���J�h���˷�	r�rX�z9���5B��u/��j�Ot~eV��p<���j*yO�]�(;���@
�e(d�u�a�7pz�A5;ϸrbT{͢'��h�匇4񔓳��?,��/����k�E3y��W����U#U=��R���s3H�b�>PM��ރ�gn�g1��1�񛷜UdE{������D(���71L�< �!�'�i[&na��Ƚ�ψ�T��Ho�#�g/M/|P�èQm�����]A����D�y��dѓ��k|=3}�9������OHdlږ��?�;0��ѼJ��g�'|�����}�T��wPb�ymeN�Nr���tJ��we[�#'t�Z�R1�PQ�gM+Oak%=��x:LY�e^H�� �W�'h��%����T?�����c��k���%��n�]�_i1i�˨wQ!9"��l
�l��a��GY�_��;�?�m9��%���?Jn�f�:M���;N���m)��r�d�w�Ɓ3��Y��ƿ�����Z1z�!�ǫ�3ఢJ=3ݱM������:���
��Zq��Dy	�����n������y�l�o*h� RqD�/̈́�-�Yf�W���zX�������
7��o������S���B�8�l��/�����Z��n=}u(�b<\P����b�-"�s1-p����{�'J�Q���G9�� ���Af+�$�SGU��Sg��v����ϦSS?���|5�#D���~�IӊG�В~���	D����TՂsB`��i�:�'��i\�
{�M&�tGX��.ޒ%/�@��i̇=�g:�u�m��8��\x�b;�ꔤV�sy1cA�Dza.7fŏ���]��􀦨i!T��Q�5�YZu7�5�^=mA�YZ������Z����0=�BB�y�$���/�k�*��UygE����:(7���rO��ؠ�`�s�Y�0�D����?�
ǣ��[�������� �ݶK��$�u۹��}���Ǘ�ū���NY�����������Ŋ��4Pt�GH-ۇG�G-ɭ���8��ml�&���U��h�?���xύ$��z\c�=��ኙ!�!(�p4	�^�n9b#q�g��f+��^	�F)�Q�dו��rc�X�/�����S��U���iO����8�'~74��ۓ$�rO��S�b�G���)o���6���W�ܬϮߡ^�t�@K��O�<%]�kT������Ml�����)	B��Xx�Xy�b4z�PaGhp�)���P�rʗ�1�U	j1U)��8�{����k�Esj�] Y59��I땕k����k�l�^�S�dH��)S��~��a��Z<^셡9��75Pw���%&��1!UN�ctx�+�c'3;�F���܁�ʒ��S�·V�>�aƫ4Q퍝�*��6E|/IF)�����@��?�٦���K�ca�����FM���aXYi��Q�����<�}�ln��۠�c�R�3���}[X]M��6W����Zǅ�:�4�/ZNj���9\�Oc����^��Pq�?*!x�P���?�Nې\�2�_@����\T<�e�v:�)ap��h�ދ(�������J��+���9<��h��,�&|�>ߡ����t�Kg���J1�\q��da���v�C�fˮL*J	@j~����6�j�W�acI�u�_/1:/[h�$���h�3�fbHN�|ow�#�_��*&f��wp�Ȃa�U]�
�Ro��#:P��׎�Xf�E�=;�d���mAwI���c)w4Y�j8�m�[��n��I%�$�4px�%P��4z�[�
Y��u��q`L����{ �D;�`�}(#c����y�O���ը�d��@�J��eL߫=�~գ����7�d�Ama��(�Uk��[�� �|}@����ox!��5J1�x��� �`�;Ƴ/�������q���-�4��zUK�E���NL����P1D"���֓��t��.���+���vǱβ��k��c��ˍI���(F+���3��v��1����ux���*��V��g�2����4v�3�̊V�x����e[���7��W_���W�=)���]|v�V�#��y��`�/�g�e��v��	��g���:��s�'����ޠ<� M2��"FQ��a�,��c��&�(q��ǟ&�ݓY<,��e�]~8��,_k��a�OӄI��g�i,��^= 3��D6n�����z^���q��+8ޭ6wq�T֭�4(YW���,��J�hS`��1̮v����s��8F�k��v���cr�� T<E�BEm�S�v�o��pt��s�3Ǩ�r��P�8�҇�6�:��Ɵ�V2���`h���A��4�壎��x%8��~��eyʖ�����K�?
4�5����8	��G)�)�E�uY��[.�N�΢$��:�K��I�����!sS�~W�{\�G������y2 ʠT��K�)��ȗ��!� P�y��yؿ�!�"X�5�ŗ�Σ�Tz� 0���D��L/DuW\�����&���(^:��'��u0u�������/�Ʀ���X�y,e�.~�nL"s�m�˟��t
�H$Nm6b���e&z����z���HO���f������g�B�zcҾp�}�Z�����;�w�炁$ƒ>�`omIҵ�3�1>� LA	Q�_3�[ 54��@ŗK� 9e�ᬭ�V�~�!�d�?C��g� ��Kz�Ȗr)�)�H�>3�II��ߊ�6IQ`���R1;����	њ&5�2�¯����u}y�WA�ٶ���O���ї�G͓x_6���-ds��b�	g,���Ĭ�b���Ҵ��C,1w=h���_��e��Gk!�W�R������Ԭ�	OY{�=��m���B��y����n��-7$�*D$�r��`�e>P�����=V��*_�ui��1�t�o��;��2h�St��gW9��1P�m[�G�e8�U����$�Y�;���MS�o�_��o�e	���ٝ6�H6��HR�fњҏ�S�Z��ɂ��6�I�����:%�Q���Q�])�b�<H"3�"3/w<�E�t*2�,7=�&3هZ*~�ȝ���]rmIFɾ!;�vD(+�I�C�օ^3�1�7�&� ���ohU���~��4��B��I�0,-Jyr�Sg����b1ƈH�p�L^yf��f��w�V�u�tu���$��V܏�cS��UF\��<B	�%�J.��!t۹�8�a���YH���1���rg;#ZJN0�۩�ཛྷ�1��>�*C��uMs����ޓ}�I63P[=�d����Hi�]io3P�_
\ݙcͮWq�y>�	�8�d;��Y�2))�����O���6f��_ѻ5Y��w���R�V�{�]]Z;ʜ�r	rџ����.�\����D��r!S��6+����n q���p�%�z� c�Hf,�:�UAE<HZ�����[�����݌�`�F��ڥ/���-=w7yBo���L��(����^�r~(~�v���6ප��da¦��鳮E� \g��(��
Xt�Ə��N$GI7֥BZ����������I~"!�;~L�g�,�b��5�o5I_
9jz��O��V�Ov���Dp�I��'c�"<BV����Ъ�Q]ՌZ��F��"���J��mAp�����.��P���H�`�dEuG�N�?Mh:$惵h�;�Q��As�6X���n���$�Hi��/Xo�I�I��A�!
��R��*�J����40a��g�:Y�*�D��[�TN���DL����z��Bz�i�0��kQ���eo���|�;�e�#��"��/T�q!���b�����:�{��o��n�4��Q�U!�X���o����V����ǰ�b��R��CD���2��w��䘯���pJ�{�棣��ȿ�ܳ<& �^��C^@s����5|K�sc��L�h8��܂�!��Z����6M���A`���>/�����l��S~J4�Pή.�]{���^�I�j-�꧷� Ɨg�LU�������"��=D���K�%����IK�B�ۆZ.�>��8����,ek��^��v�X�ʐ�`���P�lm�\�L�u٪?��@Ҍvܝ�
�e�V�t���P�D������P������ջޯ��NlY�W���'��RW� T��{*C��A�_�;���N�8�FX���3�aH �e.�$|�*�t*{%=�ג��>Ji +���2?�ԽD�&�ןB��g��>`ffW<�Lh�	��k!d�rTѤ��H�f"�5@zK1}��<@BRDR\t�Dٴܚ<Pۣl��o	IM$f�{�,�F≯�8��.J�C=P:|\_�k޹^��+�އJWо$�a��U�5�P�otz��Za�[�e���m-X�3z��/��i��{������#qW�nՌ� 
?�+�	@�7 ������%z��H��5Ϧ��*��1�/����H�QɊ����ڬ�,��<�W	��%���)7HV��)��4h�q�t�Cg���2C������W�*!����/�=����q�.ē�)��9`�d�L_��
�	����Υ_����MO��#�#�y�U���z��u(N�������=h �"�צ���Sy�0Et�kE�,L\�w��?���-A�H�v���"S�;�yR����U��;?��]]�3�v��W<��F�XUN�f��s)��z��u�	�m=z��?h�.k�y]������E�#�r�~C��)�%j��#����ģ_П���l��\�M=�&;{�~�U˴6���aB��B�b�b"A6%���O����%���!Q7Ĝ6'�
�!3�>kc0H����~���s8��Sэ2�����jqH]F�-<,"�}ڱN��Q_� �fd
�0��u�9�x���	eO]�e�ɛ���/�bl %�-y��a�D`�=q�[����}P����~/�1�s��u���v�e���%4JW����e�-���m���L��1���iM��k8<������	`��ߑ0¢��	(��)���d}�T�9p�tO����]�,�$�tuOMG:^d5�8�O�p]#Y����8�k�y����=q�-�I;@G Z�]�{,m��t1�O��)߇G�r�M�)��[b�ƤX(N䍨G�d��=��9������8��md��Ւr�$4�i���K5 K�?��ٛQ�Ca�=��t�12:��VA~ŉO^�j�D4H]B$|�:���ۖS�i;9g���+���z��{�����^���3	��������<D�g�r���m�`?�0��E��	ӗ`M>\ ��IN�4CN��q���zLl�P�͠�2��B�Bf ��f/1P#�^AI�r��g#^��d���_+y�!�f�K>=�x(��n�Xh�C�MU��s���M�����C���.3��ӭ?C���nfE�J��V����Hd#O�R1`��yS�>av��\n����<�W hiH�ܲt��2[Om=g1Z��"����u�c(�S;�=�55�G.pq��+�9�Jc�|K�C����9�
���L�̱(E�E���UݧBf�i������;�E s���F�	u����lfT��m?����.�=6N ����O�k�{�)g��J�M!�Qڲ ���(-	�L����od�ʻ3Q˕���e��lg?��vͬ6.I�s�z�.��L�%m]�`w��M��8K�

��13�β�.F����}�ʆe��Oc��O5`��	4|�'F�9H�*��q{���m:���S�`���G[Q�](řƬ�*��u	���u��A�\=�a�,w��35O���J�؈ne���A�vS<���Yl�^������T����� ���-&�m�s"${��!��D\�������K��u��g ��!\�j�W
�BH k�*�x�b�^�T�D��?��[	t	��,�Y�𰶑c|�W�����DIr�&q�2��"�ͮ/�Z�	�FH����lս�E&YWO�����ŁI��|e\��F���+�xN�K�JvMG��]��0��ֵ��B�����tz�:Q�_4˝�Z_S�ٱL?p/�S2��t��==mhU{�:�2���vلҌ�[�ǔ���T)���0LHh��۝7Ώ�BZ�:��
mM?��<�@=�9C5ڛ��,�������Cmi\1�M�@�/bx�
��'��a���~�,��N}�%�f���Z8SX.�M��2�=����ڜ6tթ���,�H_.��, �b���,�7����<��+A5�$T���H�D��`��Ωw6`/�-|�2c{��_$�%��D: �Ӟ��ׇjp����{)���iH��Z,���������H(�3�����i�,�8��O�ؠ�FH"
�~�g�<'��%���&������i�����Ү@�$����$V�3Q��`�D��IV���{����0��$OP�}Q˵S9�Yd�"�K���V:|4��C�J�wEX�"��`�c�ӈ�J�S9$h�w�S��T��v�܏��W�]y�RA�S���9d)H"�y@���nmP/M������P��Jå�!2��[G�;8����	T}�i%�w�q�.ܻ+/[����_���f(J��u�O�/q#XT�g�	@4�bc��&�Ӱ�5�����3�vL\�u��o� 1��簺 І!s͇�T�3�7�?.�O�|J3J {��[���ćL;�
���NM0VY�C�}��HԷ%���V��=e�����,.�h"}�k�Iy�3��b�e=Q�Q;��\�m�^�;qv괄�p0�y�h�-l.�#&n#������bP���}��L�����>����~&�a�Y�������Cv��,m�kq[���{Q\�&AƖw�=�������EE98�H�� .{�I�t�\�v�	+Hb����Ё� ��#e��/����/��}JLų�93fW�� �DĜ-m]��lX!ء(��K~���j����]���Ց$�2[S�Z7���GQ��"�{i�K��)�K�&<U��Ɛ��b����s�fC�I���W�H'-1F�E4�����5T�w$A�^qs����Aq���Y�SEM�Vq����Ke�!�s�x�x#���T���n�B��B�����K&Ŷ#���R*ر-$�4p�H�c���p�~��`l9u�x�i<ݱ��ߘ��Ч�q���"(�IJ�3d��hpR�Ѳn�$�:��%�#�[�L���^r��&��O���\Ij�(�G1-��]Q�����}I:�X��]R4��*��<G��㡊����m�	����2%�����k)u7Ardo���7��ip��ãٮ���z(;sZe]j�/��qE��pX<N|�"ON{��_#�"ƫ۞�Lbt������ґ)+�D���<��D���s�/���~r�mJ�ÂOÏ-�f}��LLh��$R ��)WrEڿ�Ƽ�r�p�O�i6�5��%^����FB�H�rQ%,_T���&5n�	��Ǟ�w� R`
���z�����������{մ��Ph�Sd��_��^�"^e��"(��v��Y���Z�"�'�Rwl��Z!�ڔ��{��oe�ĺ���cmݥ}�>��$0��AP9�v�!rR�9�Jm���o�r�`�v���t�<CUe�FU�ƫ���>�ܧ8=#�+��}���Z��A˻F,YH�I͵C��b�Û=�֙��]�Bt�Kȭ�0���4`v�7P�>�,��:��r���lCۻ���n�9�eζ�'Q(�o��F׈{�0`�#�_`��=	��b���d/��k(��/����$J�[�� h=�m�"�)��;1Mv�!u���9��0�w�j_�w���{��:�NsQ�(��НZ�������k~Ņp�K�=oئv${	��,�*D�04*�Z�`�B�U������z
��8��Q�*�!���1D�~��BKZ�"�HPY���c�y�K���1K���񡠭�˨p2���û����53��[��bcO#��BM4{�ON^����*Er�� ���1i�$L��+���,��F����kf�����,�QuM�,Q��K��$�ڃO�t��t_�K�PĊ�\��4��ڴq���TXoӚ�����/E�~���$:�[�0�43 ���߭Ј�����p�'J2 @'������]0�g�ks/��y�B{�I��	w㬉(ڷ�]�a�A]4����}���J������#4�*-���$�������Q�Q E��������TTn�h��JI�2�C�����Y�Xc`Um��d���b����v��3~���n���ڴF������^�DN�,���)���|��l{��$�>Pu�X8�C �A���ha^/e�(�(+�O!
�8j�����J`���|�
!i��<HJ:��$"h��y{'��x�b���f��0�@�ݻ�]�z#�|3��*���e�?D�L�T��%}��O_�눤�/����ӊ\.f�3y>�����ط�)	�Dy�$����$҂\�a0ŵ�e��m&0�?�����o&�p�ؓ�mG��K�$V�>����[��\��~}F&g B KEYr�C���BFmt3�Ld�%�(�O���>�1ε����|���\ܨ0Է�M�N����%�mC�D�Ḟ�-7��F��V��кHI<����f\Y,��>!\�\����,\��\�?�s��Z&�¿�Z�O퓗Y���l�V��KT5[f�z��zK�w�\�2Tz��cp�j�3�:�T�͙�t��I�ꩾ���b/K�HI��r*�����=l���&.V���<�JnռE4��i���[ޛ�{v���g*�b�To�J8E�ݙ�*~�D�����Dҽ���UX�Ѹ.�d��KZ�2�u�q��Ci�qq03�,AAU��{ו.��t!,OE�bZQ� �z��30*�f[" =`s%��,aZ�S�2���~Sؐ��7�}�M�Q���f�:�d>�K+�t���"��� �{F��|;H{��u�z���y})�}g�۲����h�	v�%r����@i�����qz(��n.p���B������S�my2J���4|����cl�����&GG��~�x��='������7��ю�v�!o��^5�wr�$�in�+n��G�$g��cb�I�������e˱�D%,~���֜��!E��r���B� ��S)cu�6~W�y�,�7��g�I���.Y�V�/���e�*�I��6�]��,ط>MuPBh;�鰛��
����ґ�T	
	��7�=�f�i��W �����uq���y�E�����+�B�#�Q��ռ@��m`����#<��h��˱z��^#P|跿M14�Xg�S=���^����:��wbjkl�56��t��V�氯Еk����)
��>b�&w;����J���� ]t�<\�t��GÒx7d>R����LSFu��yjc}��/�	����/3)J��%�28e�+9��
[,���!��7�T��Ʊ�X�Jɢͧ|~]~������u�Qh0qH�����T�(��=fr��D��w��U��r�GN���y.��)��U��~P�<'�R6-���I�y�h�����~'Mc�*�P^)Jɮ&&Yғ�����P��}��L�Ƃ�.$�|�G��%
��mМz�o�b�ِ`Z��j�L�h����c�H�"��k���� ��("��ZQ��Cc��i30����I�}ϕX+�3R��o�2;OE;�f��e(c���	���gd�yrk�Ejd�u��@j4�V��y�7C�8��j�+��L������(I��3w��R��ы餸��=)���V���d��.C��?�a�V�}��+�i�L�3P�{�n��`��[S��dc�"_�9�d��|%�o����@YD>�<�PP�h?�?�)���cKƩ�$Vt���ö���C����+�=�L�1/E.�����#�G�aO�8rV$&	"܅�u6�\��wT1c���4�2.�H� .�,�k�dO�Q�`�B�l4+vXT��ǈ[	W9��dz{i.X�G�'���Б
�����d{���
�۟�hm���l3|?�3'a_&����Z�M?ҥ�j�.�>⊯�W��#:y�9#=Hw�C���
�Yz5�=�P1[�f���X6��!TY^Hl���!���I�x?����"*�GEbkODaS1JS�=�#7l�Vd���Bz�)��v0�t':Z�W`׶Θ�X�˩F�*�E����ɂ�)� 3�	�'ir��@�$#g������~j����W*HpS+���TS���xm������;hF�'L��!G�RD��>���.+�HO��
k*�9�y�>��[MK����'�؆��3�� ��|�jF��Y��	���������sM�4�,g+�iF66����}TE����|�:�yܹ�5��T7��[Z�����L��N��k�Lq�g��G�z�iU{�Z[o�o�D,��8��4τ�]y��5C�`	�lQ����8�!#���!oS�� �����tt��h&B�9=��nJR�� ���!�(�H=|�nnB5�K��J@���Ċ �̌��F�zQ�x�F��a��|$�����ϰ�5�|3�c���Wv	�#������_�PM��kfW?3~�Yy����z^�&��3��󫘠�6�u��%�O>�0�S����a�~���Q-���Ek����%񜥡h�a�����V0j���Es��3蛌�?�����r!(�uMD-������y�k�S5���Z���h�p��6�����DCэavh(Rt4���ϛeh#lѭ��������	�-Sz���B�jk"}j�sփ�an�}P�z���m��g��
����ap�y�z�]̱~l�f��Q���8I�"얌���)K�
��68�{�m5�ٯJے���7@���Yfv�ژ���{�I;�?�O6�`�W�F��h����nn����׳#�����'���3Z�_XT��n���0�yD��v+o�o�8XC����z?m�}�e�0�2'�	c�%w�/�*r�ɖ�>�)��L��Wi����C��D�17+v�s6&��T�`�F��HIY箥j�@�V�B�T-V/��\H�U�����<G҉����<���X�|�A����ؑ*�,�o�nT�܏+�Ң���yl�<�2_�C�f!e�[҅�{�{��v)�)Hy]*"�����>����(�tA�Cǎ[]p�(�����=R/�[�2�D_��_��g���k�����|/����fz�� 1���U0$'�cl({mp�s��揋��A5q.��{��û�k�H���E�*�:��s[�7eθ���$'�A���Ic�dV���ٶ��0����5^�}}ˎ����`R5�b�i��)�>)P(j�z+���ұj)�.|O���,]@�@��]�D���
�8Z�qx7�\!�����6����Я��!��0sɾ���{��C�)���F�D-C�m΋���)�uV�;S�M��z����4K)P���CUkT���\�6����s��0��c�D�^;e�A��ЩЄ�vd[���#b�;d�[� ���/ZW�YsM��H[&�B��+�� CW@�{ ���������c�z��Z!�Z�w/
0�"{��wb�+�U�����P��$��/(N�����n!�=7��wFu�/zK��L>!S�PN�1�k�{Ĺ�hK���3�B��o�C�)O �����C�V����W��_��'�J��Rrʍ��Ni���{i��LX�������%0$�Pju�(�N��:���fGޓ"��#{�S�g'��7t����s��׌7��m�Sߺ��p�N���1�1�G�����jE��R�D3�T\�;{5�XX<����Y���"7�9|��XU��Ϲ=a�� ��������}?�Y��&/p+l<`SB�|�Uًl{�G�	:��=v���W}�ӡ��/t�@���̱�:������$)�O:`�[ӚkSX�
 :,�ݹ��!٩m? �O���k�����+D�,rLJ]��
v��2���RQ��H��c��CF�Y8�C��,��K��cw��{�w�*�����*6C2�(��v��:?��Тg���Е+�,�0�N��I
�{���W~ߜ�)�cb �y���H�>LNTh��Tڃۗ�;�0|i�k�pZ^y��B7o��S?*LtDi	{���e�&wAR�{M�s����l{q�W,��^��%��]�XĮ �7�*d���:��o�k#����G��Z���57�r�{1��Q�Aa� ���X��W~�w��N�P�����E�Զ�(B���I
!t/�*���	gue��Z�MB�/'�~��
e�齺|���u�
ƴ)&u��^�H �f�H�w���h9�˲���ې�+�l@�K�;�փ�"�.Z��Ϝथ*���Mrv�6SN��Z�N��82��,� ��Vo�//�AĒ��A����ۋ��r���³�+����,���
e6�5�%�*�)l��}�2��[xC��h������0M����=�	膊����3<k�W�X+?�:�$�gV���3q��e��}��H�zZZ4�Ý2��kM��Z�~C2ϑ?2���J�G�%��oe�F��_A�����3�3��On���`G�pK5�Z�[|��N><�-��3au���.�f���Z�W㯱�؁��O�,@O@��p-O����zήѦ�ԥҴ����wh�`���3ƽK���_�!���ܫe������6�ìAK�%�<hD� ��K Y	A0$�in@UDh��:�[���R�D$����1ӫ�z�!��pЛ���	�(h����Fl�%��vt����}�F��@�͇�9��˩����Ac��2>�W�}#-(��q[<M�Ru&�-욷ʂbb��B]��A�������%˭�c4��Nd�^�����<�v3��?dN�|Z�82�i�YS�!fy]�c�,�¬���%�yx&���>x&�z�X�-K�� &����:W�X�6����Fijms�g]��g���z�z{X]ݹ
�=�2jit}v����z*�LD!ΜNAD��ĬY�nǽuyq��*�F�LPZ�,�� J��"����qeH|<^��4c>�&�,UX��C�E�_`?�+j9�B����:���?��p����j� e�Ep���
��Э	�a��f6� 8EU���m9dXF�:�
Y`��N��5����Ul�;qx��E�����(��\Y�ƪ��y2�N�]�)Q�A�kb�8c�M�=�,AeT�r�`�F0�J|g�q/�dt{fȡ�	j+Ɨ�OPN=���h�^5�r]fr�%N�J��(_I�׀��u�CT>pf�O���?m���O�,L�:����� U	�֫�s�������ܮroV�~���[���@���7���}�3&�O7�p|��F���)�G7ȣTw�-^�+h�=��|4�VI�r׍gA $	��niei,��I��V�0��VO���~:�ai��n׮a�]���}��W�1�f�ڥ1Ӿ^�+��3b.%���L=����{�$� ����ڊf9��������\E���Q�O�?6aǃ�*+Gu���
�m���py\c?eK���=1�3B?��p`0�$KX��'f�S1�{f��<C��W �bNx+v��F����~��I�ŵL����x�r�݃�jW"��C�������y����������O��>]�j�9<횁��#ޣ�M�T���@Tp]�:�[�I�$+���\¾Zu9�QGjK�pEh�@�k�ˤnF�PbM<�˻�X_�0�b[��w���QZV�m'�c��P�����i8%�Hk��Q&|�	 C�-e��pu�	�ֲ5�������@��8)i�R�0$�r�N��A/ ��?8�JYL�p�{m�vN8K�Ѧ�k�ʿl����#�B��%r�7YG�bW�5˺�I��b���vA&��_e�2���ͷ��@�ڷ�o5�҉`�	1إ�#���<HN
Ŏ�l�gL���-J����{�C�`g.�E�e��a�=�y�0�騏f���_�[g�w���8�w=�)A��"�J��O��<.De�\��P�f;߆���)7~d+�z���zs1��B������p"�]|M��a;-n�Mu���o?X�(��I�7��툐K�Z0��Z�|7��'���8�
��c֮fss�����[��r�:Mz�g]YVx���*���nUV��g.��S�%�?�A���£T��!��9k0��A,��N�y�n����*G�5���QpP;�(j�8���Q��$t�e:�ku�8pW�v��\+o���E��n��v-!F[�r��7>M���)�#9!�d�N%4Su����jO�G|M��Y0U-�րߗ���<2���<�W���+g�J9ie��y����Q*��\58�h�(���/�'*���	�G�R�Ÿ<��/�8_������Lj��^��Zޖ]*��P�^��}h�,��׏}ȵ+�dW?!t�<6���'{"�ZGJ�v|aK��+u��am��<��bi��dἷ��,� �?��?��&�|?�~E�i��m��fkZ��a#+&��������d��K6B��8����<�>~�����'���}zM�H��b�7��?&H�|�F�Z�4�2����oA��c,T�[�$[�0s�Pۦ2�h���n6�[F��Tg��$7a5<����*q�����о1�T�f��v��6lR��8�ޜ��4���[
#�k!�Q��]���T�d��B����%��R}�ؗ�k�/�7;R��C*g��V�m#BM��^�t0��0��!:�R�M9�i������ �"�q�nW5g (���#���_�mD^�<�>�H����4
8G��}��t�Ya�R`��G,����=��"�
X6�ᡄj�b��O�n<�U�~��5�L�W�JZ~��T��?�Iq'�Or��H}�qD�V+�F��SΆ��/�L�-3�������C<AkQ� �x��2uz��7�����4�P=��+A$%����Ӳ��$��,/� �S[��R��*53���a������|��#c�22s��߅Pa<�2_��.��b�r�Cs�����%R���H&R��
�L�C�D�?1.��ȗ����/��>���6��`N����|F$�{�Q X*����6� ���a�W�) O��o�^*��	�@��ܓ��̃���Nӷ���-*��/�\uTıv,|<����6�y�e1�E�����)&M��d�;�=�xɉ��A��<�����0,
S���S��2����k��w��W32}�6_qy�2�8�(��j!R<���ל6�_�����@К�
ˊ(�LE����/Xފ�r�!6�'~��"��v���tV<�8���Y���JU�*ZF���DBf���hmz�ߋ�W�Taq�����2�=&8)�%T
	h��_���D�&n	� �����t��@�|B������C��E.�'c"��:�"b7��1�P��4:�K�"�����O���)Ue���[!j�A�ϓ_�}s����gz��9߶�:������:�Z�T��h���v�>���a����ފ��q��aR��c
���JUZR~&P�FM�B^�C������Ё��>��T)U�d�
T�QH���*p���)u�iq�3� ���g��n@jOŹ"�%�jȠ�]B5\�1�}c��v^��H��3���HWU�F ﲴ�%��T?���'�_@�ç�h�JM�Ŋg\��9�W���4T��}��heI�7g8w�M���\e2�� `��`BO���v�ae��o�c��ۓf��^��`�L�v 8�5�Z������1�������*t�&H&���͡gS��ˣ�΃_������_�B���<�Dm�x��� �V�b.a�E��a��f�n�Gg�%UP^��	t�k�ǜ�u$��h	��<|��|�$J��B�|;�{�r�+�VY�8���A,�Q���Bf�cH�3:x��8ߙH�gOA-!#Am囷X ���U,�fu��72��K��>V}b��
I�jd��C=�@����W�֏��j���Q�j���<"��m���,���9v�(
N��U�0_)�q�LQ�m�㶘7�����o
.�\����i]#�#=\zum����r�T��h��&��@?�ϩy�WC�Kfw��'��V�F����m6��Զ�I�T%I�r(�[�e�Ӿ�Lp޾T�����n{q2ߪt�×�xGdQ��ne9EN��(�!S����=q`���؍fb�{$m����G~��Y�4�����h��ir֋�9�*m�r"V8�Rm=����i8j�a�	ؚO;?��{;���y"Ō�}�	�T�*��J����Lŷ�,Bڛ�k��H����_�'65�"5�Yf�Z�����G6�.�P���M��l��5pz������)�@����D�Ұ�!�evj��յ�����6]O��B4��@b��'/~Ա?��������;����@�z@v��x]�ߐ�v�f��ֲ`�k���� �����5A��+}aA��#���:������7�̮zK�o��qG.ڽU�Ç�;K4C�,zE��w�_S;�ώ��B�b��׺���%ǥ[L�,��_�y��{��B�s�Β�"I9E?A������/y�rQr��F���."�3SF��U/5c㥗�&W	���5���6f���O�	ߔ~����a��L�x��?!���aGn ���I	�k&v����V�
$��-�M�M�2�;�x�/��f�?T�㷔�ȹ�Z�k�d�!j [U�2�P��4���-i4-x��[�<�Q�Ԕu��Q���͘�i��RvV�kt9�s�j��S7	Lj�>d}U�4#G![Q>���(�@��+����;�&�T�`�_s���Ӹ���*���;u�.�������C>�h����X]!����f��+�AGK�s.�	O	a3m�Q�DNZ5���K��2Ȋ�Е �5�"�)�=�By�׫�{��zՀ�66��X:	b�N��?Ń0����GHI�2�h����ADM*R�
�t�xMm|��	P�Id�4u1��#j�^�{E&�ɫ[��gdWX��{<��c�g��M�g����g�V�����h�-4�N���c����i��9�4�;�l&ېN�Θ�Aot���@(�ݠ?2��T���a�ۡ�ԗ�&rsZB��Y����O=p��o}W�����6m0�TAoZ':��g��>�(]Q�9�������bi�V�S�L_�剈����r��C/l'�EP��@tҜ�r��$���&�/0W\u�z����$.���@䉷��$�'D�jI]�8ϒji9F��\ç$�f�*`��v?9r.	͖C�V���mP���V�|���(�V	�vy���5�&�����'+�����l������r���3��f��}���H?�A�C5X�AJx��a�5���$K�z��癋�
N��n�	�_�S�
���kou����Ր�T�e�{�6%��R��I�!]ʀ�qbe2/��p�*l���l<Dq��[��,�n�ԄS������Q��!>�^��į�%m��P��8H5|�E�C���@Gx����	�9��zb+���D� �b�1�g�1d�>�VaOӄLA4�kH2�����Oi��� ������)��Lt����̀��`@��.��&�G88�,}�pɿ�6
��>zi7$������.ɸf�YS)Ό���w�}�����Bg!�dk����� �g���,cv�9�����/����8��3W
�Y����+�:s�4�yq����Eb��Q^������$&�"g�c1�H�;O�y�9����x���B `߼�gO�!��'�{�g.�&�ϐ��;�.��� �ݞ#��W(��X#[���f&�����]���d�1�h�a�Κ`�����jWI�}0z�B�eϿ�0z��ʿ�+Ia����:�Ӝ�#<�w��U�t�Tߚ(a/K~�
�̋��ƕ������07!�*"�Q\��,-�m݁����놿���]7���ɩ�qy�p;<c����/�&	�f���Z���4��3z	�&H�^t4��6����2��9��y�J��N��y�>��.~ݥ�Z)��䨹g�~{S�WZ�b�䜸^2�|��ɦ�:�vH��$AѵBI�#ӳ;C%隡s�a��$e��V0?�Di�Y~#�����[e������>�*R!x?�Kɫ��~� ���^Es�G���`:�]��M�C��5@+(@ߞ����d�m(BhDA��1�D����32�溑)Ȥ#2��  *��$����	wv�u���$6'��$o�oٖM�ys�3��R ZP��ݼ�O(J�(_j��H��ZM2&����Jc�t��T��Jé�A���G����}O1[�~��D�����&Nܕ��r[ _+�i��o�U֪b�f�Q���A��Ih��G�U1(dMo5rS!s�����{n15Յl
[�]<J����˛�ئ��l �_-O�����eT0g�J@'6���bI��5���$��+���͂N;��h�d�ݝ��|�$�3 nF(qV�2U�g�e��3����*n�Kf�d����2mC��)�2+BG,8Q�)�{�HJ��Q��f�NHs���3��3d��1ty9	����|��߆J��n���Wk���xY���A���uo�n��'���$�^U�I*����)�Y��J|���];���c�)[��z�L��0W�ѱ��d�(!�{{�ks�307U^�]���!N}1�hR?��H�ފ��Z�Ǝ�������k�����j��_���V�9�v�����*�y�71kp��/\R�6W�~�"8��/���q.��bJ�j��В�vVk�ݮ�n�0�N��z��'���4��?P��1�y��X[��_�*Ub}������2�v�K�9��_��5�#,Q�(��~a�f.N�8��}��*
z��JU�:���l���㜈���lD�zatt^�-��ʴ��Q�?�.�����\����c���?e"�U>�I�6q���׌�\�R�%C!�`��4�[��9�{��v>[�M����i�EtT�.;9eP��~�Co��`V*��Y�F�?!)�Q{�&��喍�v�ڇB擕-W}!:�GP�ߢ4�����t�Fqw�d|�_�p��<�c�v�%�is���J�=m�"6�Fk�Bx���R�ihE5usЛGWF�UO��TbB��d1p+���TBq]N�W�̣0�Q��ɸh%p�d�tf���G��:Aup:)K3�A��Ugv����/�����$y�@���-�<�'3��=�v^	>.V�ۡC`W��_����������~��ᗢ��ld�H�aYM�]�N���㠫�K���-Ж�4 
x:��gr��,OWl.�1}G�,�)�=�2�DcTn{zj�����us�.I�����HI�bk���ӢF��R��ޗo�T)�k����۠�����a+�, ���ps=9��^c>��L�n2���^����@r�k< ��N���&�%�G�f���e�OIǁ�ӶҪ���Ȃ ^! t�����;��Ҭ�P��#�S���;�6?��'j�K�����1����/�|	yo�e�3/��#����e��|�T�����Q<je	[�ئ&�Ek��C3A�.��_zǜ�#�V�}�<ZDK�q�fItj�P���D+�%��W��p�e<Zb��훰��MTA��>�ޘ�����~��l�逺��j�:�s��7�퐠aB��N�^�(9�V�Ipa���Py�)>����AP��;·��A��$(1<���D�ĢH���٠#{�ތ�����ԏ��ɪ�Ш%�����LתX��Vbr�9r����f�so����e?�'��>��_��i�<(x��~���a3�\H���ᢨ�K���B��F�ں\l�%C���˸MC�Ȍv�ׅrO��rx��W�s��ZJ�{��T����<������Ah���{Qd���`2q5�U��D`�>�/ႀ�{f������!L�����Z���⁫��^���O��&,_�T�B׋<��c����Ym�;�2vU��3wo�%� W)��~�q��U%)��8��K6_�E4 Ab?K� T�uT�7��p�<�P�ĝ�����~ &��σ
���Ճ+*Qw�U���Je���Y���2�>^j.��ze��.ܠ���K�(��ܗ����1z�J"��,�Nc��\��07���Ec͔��$ޜ�ȓ��R���{Aq�
��)F�0MA�K̠9Ug|x~�� ��Q��5.q	����U.� ��ࢄY�4b��XH&�Qg%�2�3�JW^bc�ӟ��@[�\�0tmW6$�b������c�Uzz�m�,� (�Oq��c�k��d����5^�����ו��*�2�Wj �b��"6��OWr����S�V��N�U]��C���tΒ�]R��h�u!�����l���4�U�@��}3H�ք� Ω|B�{f��~l��&��fߙ&^�e�͸�O��$g�����Cc?�]�k�^�y�6(�5!t"x�&�R�y�/7d/h�ĳhX�A%���� }��JVdU�o�Ѐ>^
K�Q���	��� ���u/WEO�s�C�^��ʿ\\u��s<�xz~�0�>��ф?��P���޶�]��z|%i&F�;؟�VS�����
`�Q���||t��]�a��0��K�T�;�6농��&8�3�|�0T��"2V�l��~:XӶՍ���^���z-'GlW:��/��|C�+E��W�U�Nm�����4�vP���
 &Ph6t�1g�ZGm^�0���^W����Mгr���Z���2�~&��D�F:4�4�z�� ������z�c�	�^M��`'52w�<$ǈ68~�)e��aP���UxiDీ��"��9�؆�«���r;��j)n5�+en�>m�XtN��g�큰�.�+����E75nut�Q��}���f%��=#�Ր� ���^P�+F(C�/%�e��
И��3���}~_wr~m�	~c,��-�%텤�%"�<'��P��
�7G��-�'��=�B�8���6�hգaq����;P���v���'��:u���������GŹֳ�������y�U%P�C0��@��sS�D�D������V~!H��i�+�E ��(��a2/�����������54Z~�f<����!^��X����7���oQ�����d��Qtɪ���5�%5�a���y��d��wf���c;ߪ4��φMQ�
a�u���2�A�_���i�5���yr��@��ؕo��<�>� 㖱�V�=nZm��/N�+��jP�c2�������/��q��1�2x���Z����h�UV8���s$5�W� f �#f�j�ɨ4Od�^����&LXѸ��������T<9V��-��~��!��â�w/�2�
������5��h�Ĕt�΂����,� �x����.���~��jjh|O])��ZG�D�@�k�}Ť{���gR�&ӗ�B_�0���01vg+���E�����G���<�����]t׸���Ev���*�,�I~�w𼶨dWΘu�G8x;�y�V�bvp�Kш��m�ekF/{i��Ђ� ۖ��5�
V��k!��J<3��:����H�H�_����,���gcqA7�g� B����b�?`&�D����a�:Q��z0�qiF*��ū���_�&���*yE�1#����D	#�4�,�kf�e+��W2����-E Z��F��Z�|h$�Z�����R���N��?�6/F�y�/A��s�5Wp�P�@*4����@������g�B?���深��;�6h3	�P-@�l�-��ޕ�?�l*<��@�Z�	��w�K� ����G�Iy�H-����l~�I֮6�A ����8_��'��[8Bऋf<U���v+*	"�;��J*-�aG��,��e����xa7qAqQB�i@cGA/�
�un� CjP���K�L�{RH�ӟO+ggN�:�x'N&�ky�fd�awn�Oڊ)�3�r�@v�f� ���vm%�X�ח���CCCc�lC���hXk�D��G?-�5՞��}�
[�3N��̇��o#J��`��{,~�m6�S�O/rL�ل��_�O�Ϛ�;
z8�g�Q������:Nf*�vBaQ�q�'+my�Royv#*��9.&�)���G��?�5�%�0��fܟl���%t{yr��6j3�V!HI��W�ɑu���'�*7>7�5�!s�M��3	�$���󜅬�n��
A�0+���7�G�����~��d8���"����`����o��?2�<�Bl�"�l�8���ܓ�KZec��Ķ�3��~��8���t��!v� �K��H5
������UF���C( -z�;�gsɴ�|e��-�%��TȚ5�T,tc��\U^�w�G:M� �Y<ID�c�	�P[n30ќ��P�l�T:JS�7o���q4���j�S~^zט�MbVڎ)C����'kp�ltW}����ɶ�b�]ʔ���U���2��)Ws��fLҬ�%�^/��_;�Tt��1H���cUFv��,4s��.���bFHO�t�2�S�[1��3�0c�Z���$ C��o0\Z pay3y��5��J�bĸ٬QoLǝa}K������*��$u	�9�PH���z�s��n���� �~"k�JN�7�ջ�m]d�9�AW��������+O�C�a�!B3��0XX)�)�3�K�����cދg�3jcjeС� �[���W�o#;��/��,'X��$�\1gCK�D��Yx��0|����S%�yh��"�PQ���Ne~�G����j�����Z�������669p�~��k��vZJ�i��{�����Qx��i��ۺ��T��s=z�}OF|���=j 6��~��\��30�!!.'�e�9e��+V�vC�x�-����0�d�pO�eT�V��B߯hn��n�Ŝ�e8��'gD��/�Sג�'��B�.������lт � �?���g����%���"f����������G�2��6����+���J��ʓ�'�=��8~��?�a��� c��p�˙��U�LW��$��v�<8�nW�p�U����}�
,�kT�f�HQ��Q<#*�?�е��3F*�_=w����5��5W���ݛ�j��=%���qͫ��m	��4L���k��܅E�-���n���1����c2���WQ���]ǳ�	J,s�PV'�ķ�r��v�)���5$�<}��ֽ�,/}�?�doF�5�g��X)�ZẎW��y�Q��vX�_w#0��
J?y%��ZjQc)^�Ue18��< �y����Ao�Qև�U�v��a���4����`�
^[������r��MZ!mș5ϩ��dO�h�� l�Px#�p^7��m�0cј�~g�"��������aҜ���ߓ�*pt�_�x�fj�X�iӸ�d�l������7��M����H�n.^}��� �l�SQqD�F�`D�,��_�晹-e�����I����Ksa�М�_�p^b�נ�by�n���*�^�n��^0���� BG����9C�F�S�[�2���>�@P�4d5*v[^��:v���a��m��:Y��j$\��֥�{�E���z�����?�rC��Q�'��L¤��ytv'ŝO���4�[�X�=Kj٠�.�*�I�����3�g�<��ۢN���(�Ya�U��P�Zy�q���OJ����7���=Z�0&d�f%~�0*�/�em�o`~%C��$69+>�)-�1��n���x�v[�󘓡XU6?ϻ�0d��3��?j�󁵉{�M�$����t��㝸�':%��C�bx���#�D��[\�	��pF���e��h4�"CL��R����SvNv)ڙj1���(��e�oH��dU����
��dX��v"��B�0e�(���w��>\f.{M���DN�+�lS֭���L��] ٳ��).��g %�s������XܕxLd����Ŵ:�|�)�Hp8b)DZ*��7q��}�J^�a�&OW�M\#��c�V����v�($Y��tl/��Z?G!A�6zQ��Ѣ��$�ښ��0����x�&�����r��y
R���ᝇ�L��P��"��)�����7�?:���1�9?�7%�0S�J�A(���L�3@��;tHI�8Dc�[&B���J�5��D�ԝ�bk���|'+MB��r�6I�[��pn5ci-��	����͂!װ+���B`��cꈝ����G�U�W5���uΝjy�CU>X`���;#�aq��DUC�����ؾJZ]�-_�{l�m�<9�[H��/��(�~���g��H�����b�����p�o�W��HB��;2�h#���w
��ϱ���G*u^-��#�u�'4&ի����IZ���D֠�����W�}���,�R����1�+��#��QmȤ�U�E�h p���Z]0_6��}V�>���7�����̏%>_q\��(k7�\��1��t�a��<g��P���5��N���A�ck��<��-������F4�(�a�$�g;A��/���K��k	��K��,�r��A�R�l�+�n�� �s��ۿ�%�����:�9S������ؖq������	��O��p���:&��_T?���x�32>Ha�D�+��K|aXt��)b~إ���$y�k��̤��r�;�yѳ�>����o�Z�*1ı1}�aass�GWp���=RFd��K�㒗!�[yK�<���<�pj�aƾ9C{��z�0'O\!
�q���zL�-h���Fzu:��OciМG��j�c%��v�,X*��yuO&=]�(M�&ת�YP�?��*Q93{�?Ag�TH�]⽅���]�-P��x�p�a�&d�׼�@\�Z�SH��,@P%|�~Q	M>�$f�g�h6���%p�0y5y�NY�h�Q�W�=Yn�=��E{)�Lvۭ��8���F�F�#m�xIb@d^� l���f{�[ ��ʺ�9+�&�Kؠ�عSiP�\A�Ŭ7��62�NlX<1��0�.����@#[-8]��Y:;��A
�^Vp����ˏ��[뾤�MP����4aCr����c%RT?�]�\fs�弶�q�}n+iҵ��G3
�����G��O@�oZ�dA֭��������(h^j�3��)ҡ��aC��(�	o��8N��0�GLA��m�>̯w���(�؅	�β�چ��Ƕ{"J��#J���&��;��}L0N�#���j~nTg�VA�����}0�e/g8Y�M�L��'-�_�ˏp�E`pR�o?�M吐����������Wu�%�Q���%��ב`ʵ��h�� �'`�|W��4�bxX���j� ~V%<���o����F�E��@d=��*a�w����s�:X%ߺ���}ѩ���e'�w��5�T��(��q�3�mGj�Z����-,���Π����k&�:ٖ�,8/��}�>�AϨo�V�)����-@����~�R�/�8��t�Ԯ���T���o�d�T9&�mmO�F�o[���p˕���	.��?����[[x�����y-e֔9��e����*M.��H�rۨE{��2n3�x�Q�V��K��ig[)�e�?9�����+�6��H[����L��&��>٘5��%� Jb3u5=/\����>/�[�������b�'��uf�#���}���2��㬓ai3��s͜)o��	�4���i��z�`kH�UB�Q����z���x���Xe�W�����yAX��9�xa��H�JO+&�Џ�h��Ah�u��_EnU!��J
L�4,nn��2�;~�I���pf�;Z~Y�Ǜ���'��s9�l�:4�kK��Qq�- ���&w=����M�a�V�tz� ��.ǽX;4h	�B�U�H2���x����2�j�*���w�$�� 6��/^O-z�c#�0��p��$�r?�q��"-���|�;��5$�G=զ�}�$[	sM��yeHc�d�Q�"��"���,�����F{��IܟJ7�zo�͞��N勚�M>6�������E�\��`���gP��^�� �v����4:}=�-�A�~	�ʓ� ��-5�w���=�	vTa�V��-��3|�J(?�b6�-hj��� ̢�	���v_��]���o\�m�]Tv!BXNlƕ�������r��\�`8%~�:���Q�CA�Dd�\���v�s�KO<h���%>ժ��&�(m~��]�O$_A2�v�
��ϗ(A��<Q���QDi���e�������b�z�dه�����k���E�𩧙���2;���E:��&2���\V/\p ;�N�+��V�Qw���ƿR(����@\�X��Z���\ӮvM�H��!ZP�6:Iwj ����#w�ۆ`]V��69�_�g�g��1s���IR�K)������9����-�9r}���I����*��Mv'�G2|d�'�2��3��ٲ�3�i�m�-���@����WJ7�]+o�V�[�KU��O��
�f�l�`����dƓ����j]ې�?����o��1wc(���� �]j�"j�R6'=I�Ք����h�E5��F;�9o-��M��U������/O( 6.N'���7���=j�r�sBa��1�
0D[!��*ʜl�Op��m ��>�<'�ڱ��9�1ݮ�!����I���%nKE��}�����3HӤ�8��ͱ������-�<�xA�]��<m2`��I,������|}��CM-��i+�PJ�و�Z�?��K7-"��Q�M�5,���SU�4j����]���C.�&j��g��7���	o�荪RZ|���=�Q�@�暘�Y �����1	�S�f��ٟ�M&��u-o��Jr�{z߬d����q��_��p�_��f��DA+�5 Sh�?��V�L*L"�G?� ��,��݇g[�K�IXOZ7ȋ��' i�0����汔�Y��~,��`K3
�����0U�T�&: [v�[��ۣ�̉m��_z����#�8)/��ɞ_��4tG[=��8*2���C����L��[�c�<~�I�J��0��X츽���3����-����,��?��MK�������l�E�~�:�g�����k4r��3����)-h'b��Pm�*	T���UnW�E1�$�-�I�<L^9p�k��/)�'�r�Gq�D��л�}3L;T����'�"R'�7��Ы��S�f�Fe�m���U*����y�邈3j}�����zxX"XB�>�$�"x���Hjp���Mgr-���Cb�u��j�\��J?�鯓G9�NKr8pW{�*�?]��p� �C� "��&Xx�!U<`�W��4#�l+X�p �Ty��8���X^�f�a�nf�K��K=��>�ɪ�o�L�H���O#����d]Y4��f��H��dw���u�kV���x1 A�eݸ�'{��� گM �!����l������u��P?w�{,�ߤIf͗�1�����D�XLPK�&�\".ۥ��|}����'^���⸮��|{�,������z֙��]�J�Q�yΫ1���gJ]�	���k�=Cni)��[l#i�p4��Uo�O�1�	��k�{�fE `��T���K�f�LB�oð�;S������a]�V �z�����֞v. �Q>���p��-'${�������<�Vɮ���YO7�?�M�t@ ��kO�Kp�23G�M仰�u��M����I��u�;��g��*�X�n-��Z�`^gN� a-��j���v��-k�>�R��0H��}0�����؉�C¬p�093,ұ�?�~�zʾg�\�����������Q3���-p��Eza������>tO�J*�ou�M<��G��u��/-�j���;*H1�{*:�:�h��[�&���-w������&2�w$���H?�
��7ҭ��������_	g�
�Ʉ��׾�WՋ7��!xx�qj���},`+�f�J��*��k�^�/�)]M�Q�?��j�M��)E�a��b�Y�)�iv�{���Uk�%'�ٟ��ǂ�դuۇ��L/eH�<�Dگz�����瘌2X�jor�.�s⍥T���d[��aZԚ;y���2>9�S���e��-MbV%W~U ��p4�?	�6�97W�:5S���	XyZ?�͉t�X�>	�AU���`X隍�O��t����$�;���Jyl�Y+�GՒ0�*s�(�5�S�۶D�N��wp6�>���0������	X�*)=�z�?eٱ�%�䜥i�?�`��кߤ`+<��.e�,k�o+�?GTF�����k2ɲf� 6�j��zo����u�8x�=01�m�����w��[�=̀�}Ŧ�?�"p5c���=�����$�,��S5Ą�y��MQ/C�6�������>��L�ڈ�1��Uy2�B�-������*,|�eh��MI����zp���Î$4�ѣ��_������6���d���t� ��x�R�hd,�,��4d�Y?��*����I�$���4���H�ĶХ�`���F���G�B+�v:A{`�#*6SD��{%���d����D)��
����1���M#��I�)8��èv(���(��@��1��ę�L�-�7L����~�`���G�/��/&���ۯ�ZJX����ܭE�&�:r��%�ù���1���&/s] zMM��Q�up�RqFbU+��Gh�U�Prm��@Es�Fk.((�=̼��!a��ԸX����CHX�$,XO�$8��"ײK�Vu�97?���K�D���m��/��|L��P�OL9uFVȇy�q��Ɯ������^�M�W�V_ſ7�ǵ��
�����Z�\�P�Y���Ղ���nAa7A����B�Dٳr�7�) �_S���Ͻ �3z�D?�EY^R���Y&F�,N��x��~�	=x�ǻ��7�F;X�\5��lv^�����1��0��L?������k�-E�� �F	��SǜhE5�%4����~�Z���sy�|\�%�4�Ǚg&K}%f��|��fjw9Wu��d;��3<��ڥ���ǓMT-<T��H��u�FN�ߴ�xw�k�X��e(�b��hm舮�Xd^��6"�T�1V��[f�R�l�?3�͚����<V�\P_����w}�uyy)Yq"��wYJz[r�$i��N�K�/�F������S�Z\k�2�D�{�����n):�&+�\�E֙�'��K�H5l8�%���S��I3"�o���_�}��K����p����� �񩿸@M�҅��f~WW~y?���$��w���NU����q,l��i+�-��Ic���|�&'�h,�p!M˅�fMA@W�w�"��x����㚯h4��@]2{}�v��W�} #����t�Ɲ����oY��tz���:�d�"Ql�1�5 3�4��M�����'���H8�(?�|��OtS�^R��H��t���DWݳY�Қ��G�Fq'��F�:<�7ņ�e�+m�����<����"���Q����QԢ�뒝+�r�B6v� �a��Ӊ՘��1��Rs���2O��b|���្����9��^(�T����5(@S�!�{`;�w�����p�"S�oa?��hÛ�1�^�%*�-�~	f�Q�`+�y�>�7�{j-����ۗ�9es �Ha�-Q���w�����;l���+�(���K/�PK�@h���vSt}���5Bx!�����ѠwmjF�e�Q�@4X�T�7��2�.��'~��Z쩖k��ԭSp�>A�9
�_�=�$ߋs[
���Q��=����a�n@�To�Jb�ܔ�4S$kj ��ƥ��� *T�3-�f����a�`�Xp ��7�i��L@��R&��E��J���E)�h�q�1G��sE�Md99�iy[�4%�5~�:���]V&���&9'l{ř�KaSue����InM�3�%~��C#���f���8����h�˺��X�y�|%���Ǥ\g��+WݥܵRoͤW��il��Nƽ���Z�B�o�3��� ��%F�J35Gʓ@�i����+��������_M��"aŷ�Y��R��<�i^��]pE5�F()���Fʞ9<b5�_qF������|�� se��o��`�/1M�q��g��躋Ʉ����],�m����o����3�~tIA(~w�D�B�n;�e�D���<���ɐ�-g�R����A�BjN��/�������A;�8J�:knlrH�&C~�	��ø&����ׅs�� �8���>ĩ���Z>D�D(�w�DY�_k[x�Ӹr�D�_	�$�$�n�iG��}D�Հ��Q�Ǟ�侭=��[���4Xx�1�|��/)�s���7���,�= �!����m�M�����J�$~4���l��N�a�I���n���I���Ϸ�ki�d��'��|�%57R�� 1#�%����"FҶ�NI�q,�D�g����=�e^ �1}����eRuP�a�LV�;v��5J�2��B���y�|���m�3��P������h�޿5�'*#1OM��ҲaX�CK�%���[��������q�1H,��\x�G���5����S�F�p"F���3�6�_���i��8'"e�U�\]u�6�����B�Qf�� Ƽ���\�΀d5�x��Y�9�L�� �VSM._j�J��M��É��;[;1�+�"�O����Z�V|[��+���#Q�۱�L.�2Ȋ,�� 4؇ ���c�RHjY��(�I�o~�R���Qȫgb��q:E��0������zK�����K�I]��J����v�9�o�Q ~�CA��l�ጣ��~)}��'�桄"�uſ(L���A%�ՌaI(.v��溔4x��D]j-�I��5!x�_��y"�<�C4I�d�i>���"lc%D
�X�b2�]t	�K�>LY"	Zx���sg}���q+���7�p�{C��>Ifˋ�[����k�V�x��YO�XI*�9�r��%���K���)uQ:P%��H�"& Pg�:��^�v�֙0�D��~  M���<\s!6�<v>P�?���wY�"��H*��tb*!`l�G�[-j\"��Ϫ��
����5�6|�Y��h^S��n�����:�hM���y�;P�P�/B'%���n�g�Q�F�z%��ylH�\s������oA]'�}[PNu�꽐v�!`=O��h��|��֝�vͯ��0uN���*'�L�� @�u� U�e�ƔD�i�������� ��?���F��|=��<qz��_�M��� �0��3��=��k
�~/$���_����'7	���t�����˖k}Vh\&1��u�`�A��ujuֵV="�x:?j�G��˹���_t�ڡ���H5�1
�)�TPK�h.��!��v�$�+<�p�̼Q��F��[m^]�4K��2��D����#}�*K��gt�Y��D9�O>I����D,��\�Y�f���_4꽠�����a�� ��]�7v���@�E�fv mGD����� �_�ˬ �2 ]��C�l�w.Ƶ�������]0�L�~�����׊9ws����U4^h�A�ur���\+]����gkI�U!)�K9l�r2=_Z/�yZ�f��)<V(̀��h@�īT����:5�v��S������7�F��;��sC��cϡ��[FO�6�ܔ�^鴄R�H�H| �ŵ1�����8r���qO�擰xf��0�\�Nz�6aw%�_���gX#
�k��V����`>bXV'�5��ƅ=��/Vpt�:A��`N�;�Q��}Wܛ���"i�y�U��;<k�3,H����ںj�� �r7�)%�������_tK��hr�f��d*#�?,١��Lހ��U`�E~A)�Ó���7�/֣z�O">�
�3\f�n,y(��LѨ��q�4�Ý�O���x�u�_�
��p�S�%�寨�?�]^:��f�x�O.�D�yB@:��X�pu���t�ϫk�ѫ{*�z�&��������m��#�j�4���� NW�;�[;�
<F����1C�	v�H��32�*�x�̗�M<�O�čq�(7�7gy\��R���T�U5Khɂ�^|��w�8�l�˴��bGpK�)�*<�I}��'�W�y,ءJ����)7!�d��Gy9��-��<,�fJSx�Z{�x{�<��څv5dխF`]1$��@yq�)�`0�u/�������ҍ��΂g��:4 ,��ߔ;�7�;n�W�=y�Ah�Y
"��=��� `\^a@���L#��ۧ>Vk:���2�B\i�im�����)����������@���*�4�I2��=�����Ԃ�����Fs�Ʌ��r��a3�����Ȁf��k�3*����+�*�nA/l
4���J���%�̑�4�� ���uE�1��;��t��V�VR���3�v?Qo�v��OpT�Q�cog�Zv댢�. ����e�Z���/��U9WvSmxA 4���aD��װ��+�C^���)�=K�4n��.�x�=�]��P�ܖ�uD��#�%����JT��^*h�}�M��>��J�R�*]�	�R�E����QԨR!+Xի������.��JQH����2�%m��|$�O��"_�gE�%�g�l����1���+`Ճ7ԎG��p�4�^v-����<� Sݗc`Q]ߒ��4�0�'�LYU�0��Nڈ���j�W��bC��ϯvQ͓g4�L����Ue�)�ץ� ����+RK}��������;����g\�{��IU*c����^ tΖ{��h�)��"M��}i�R�b�4+�G"���O��M��s�����g	�	�=�)�3��*��Ӱe�d.>D;������u� �l�<A�]+��p�F��Z,+<M�~9��� ��^5��{����!N6���M9���������1!��e9ƢcO��W�6_�1�UX�/�i���&���m�t&��k����1�G-#K�jr��|Ŝp0Y�R����@H2�qҸ�D��'[����? Hb����57+���]xxX�T^�;��0�c��5c^����h�[\�	�#;(m=
�~���7�BV9�
�I�]\��-r���*v��ߖ���ݵB83�	�w���B������kP�48�k���m���+���c�JE 4^�e�p�o����jf%�a�-/�Hy��W��<M����[����ؿ��xp�m��S `���9�K�r�jW��i���y�܇�ͱBϢ�L㺗�l�W�%��1x<,�t�6z�q/����9���a�4D�hKY��e�d��Ÿ�E/��^Vl(Sw��O�,�y��l��69� �J�׵��w�,<3���p���߷KA�R��O�I@���V=�01��KU���ˑ��\�ll�P��eL��ԑ�VR�O��p=��}I|Ypi��34��گ_L�L�.3 s�Wdo��������ɢ�3�`y�aØ���F�l�q�u˓A����9�G���5z}F��U ��50��A�nZ�����p��e��~�e�����+b���6�`ǹ+��\}��u�a��}�����|Vlؒc
��[��u���h�N7��PLc�R�RZ��i�Ʈ�J����D,ѽ
�PkםKp���1���(��ƕn��&�Y��NO��D�d�0J7k�9�C��ڊ��,�޸�����GfB^��j���t��@��n����cj{�z����K!���D�g��ɭ'�ThD���:d�+�h�#���y�j�(�&2���2v@2���A�J `��f�UJK�Z�Da������N�^�(��ٽ���C�>��J��$za,v�4�w>����^����%�ܛ�Y]%�Ttç�4�c�r�G��^�^�v�G�^�W��;���k���l�����������T��/�dJ�~����YNL��A�])��/�K�z!��f=��S<���b�~��~�ݴ-a�� ��A�UA���^a���5�t� ��Ll�t�r�����F
15BR��ɼ�d���T���(�l��!��6G�����
���̈���P�lr�-N�w�K$-�Yuol��'�UK�KN���ӥ���/+,�ɗ�_w�j�b��}T�n�E�1�	9h��p�z��4�c��l�@$&`R�����K(��K�7c���م��* �+��L{��^�B*,��ƪ�wFa(�X�DG������Hc�YV*e՞�[fDJ�����~��~OF"��Ul����rٶ �3GY}�"kI]��/9����:������Y���P���h�V^�F��?��ȹ~_]�*������9'a\$�t!Y迾�5��#�[
(����Rs�.s���|t]��bD�ٸht�O�-ފU��!����ZSo�G��$��N)�AX�X�� ��]�g���X����c�˨��'�!�4ʜT�ѥ�F���(%~*|������,+v��xI+c/C�g��A\I�+~%g1�,�tW��Y�9^��q�r�!������dT���������7j���D9��S�i�Z�� K�B�]��"�P`X�vXc Q��ي�4%��cUxGy��,��&��!�����K�b8����Q���9V��QC-k����ko�ZV�R��Xɳ�e~=�[�A�4K醶Q.>�V�L��=ZAm-��Uڅyz?x��S?Lz��U_�=��zL�H]��wIXP��*���e��h�>�B@��Ow������U���/���qUq�ѯ�Pծ�/7��{S�-r��+BY= (O{�W]/����.�Eu�:,���N+���Q�l�D	�q3(�7�X~{���p�Y���ɇ�Q��W� ���g}m��ݽEv��Qd�5选�M�L����9"�DX��{�@Q�U3d[Y�;0jZ�t�FCo��]����)�Oxf��mݰ΃]aj�7ذh�d��+2b}� �Gj&��Ϧ�ࣆ�}ڿҦRsG�C>�E��h5�g/��(j��/|�V�Ԍ2�N��8�|M�j��>Ӻ����Z�l�&�ʌJWA��&�ڬ8�Q��ėh�S���EW�RV=���t�֫��Mzܧ�-�+?�������ߨ��#��}���C1���7�j|{�v��X�p�L�/k�ɕp�9w
T�x���=HY��m��OWܟc=�ו�I��w3g�F��"���8�wl3Z�$�b�#�P���Lh��53i�/��%���z ��Ɛ�[V&k^�%~zj�>X��d73,��~e��N��*�M�8�	rZ:������A�R���h]���98aĳ��u��-*@�v�w�)���.x�ϫjT)�VL�n%�F�X���Y�
�̞�EEQu`I!9�M�2�p�!�Z��W�������g?��KQ5�>��%9��X%73�>L����f�*���~J�S�Э�/����\'���L���R��|�@��"���ut�X�����Bn���v�p�f_,�`��Anb��*��H�U��� R�`½�ƈ�	�P�Zv���m�U�|����Ƿ���JT�:J��v麿��BLL3�������=Ƈ]d��쐖>�a�QQ���|hYm|�!F<�����1҅�gyvM�^m�[��ن��>}�Ns/��
h/��WB���#� �=/���l&3I)�ߺ2L`W�g!D�>4��,��Dx��)`&Ǩ�ey�w��m��FT���Z�,REh8�`�5[Fx�ԡ%�q�Bx;��Y��HM)&�D���#�_�xA�ן�x����ChhՏG�U�V��*&}�4D��<�C��S| ޜ`��3�c�N�?�ui�=��8���d�L����uߞh�<��]p;�Ĥ��gO!p�X
�!��]\�'y	�C��P�,�;�A�H��C�0 $0�l��(K�*b�f!ibŴFP�sJ����pp���a��WT�)��3L4T��	�I[��B�K����	|!�`K9Tr� �l�aQ�@1��p�WWaa�D/�s��C����:��w�T�f"�Vۅ�csG�Vqa?��&r6�����e���`c�7(�9_�� ���P����Hw���c��f���Ȭ��P�3�A��#3�R��i}s�)Jxz��v�_�1�S4�`�%�>��E�1u�A��oh�MC#��+�����wd���;��x9"���CQ���n���������0Co������ü���&]I�/ٸU��hDN嗱)K�^[�	���57�W�#�i�+cQ@�[HkN���n�(.�|��o/!�zJJK�X�S�/޺��ABb����r�k���|�(*�z�H�����U���_5Vg��v���>{
����<��o/i�Ⳍ�Wh��p�|�jsru�c
���~�3 �5�O7<�]h�돤D`��x�c��S&��K([^o���9k҅(���9uN��ԁ���N��F��|���q���Ћ k�`�7��ѥ(Co�� ��Y�_�b���̻�%�R�Q���ok��my�eu˯���Z�����{@);��ɚe�:�Y�y,]6W�"�/rʠ�F��y����c�S��(xQ�YR�*��BGh�!\-��8�Zz�K������Ė����v��ƍ�'2ENH�b��B	i%���0��[$�AY��Jх��
��D�_�d�({
��4��?�;�{�F�?�h�T����6 ������;�R�8u�?�}����C�g~��0�b��M�P���|�	R�`�vQ��
�s��y>����l�O���B� ����5��]�����/I�U����q��i�@��vn1�,gX%a��Z�
}lSD`�t�i(C�?C��Л?^�0��P��b�y5�WD�7��\������4����߽�U�_L�i.�I+S+��u��G-5�@�.�MS�*�Ҩ���SDnҁ�r�f\=��Ȟ?�ȼ�NmeƼ��a����P��q �z��?��p�赍�	���Qih4����+@��SRZ�L��:ad�|-�	Z�^2���~�e�+�@�!:�����f�Ӏo�>'9��G�� 9��n<�G�H�^���Ͳ G�Y}<�� 3��M�0|��D6'>�)*iF�P�t?��yE�K�:�2��^
%����"+�{1�y��CR?f��0�0{IH"��r�Y����Dc1�ψR�
��3������*��ȹAV����d�t?�X��pͫ�$�
	'��s��0kx� � %�lB��M��W/'�������T�� ��'���z1U���
�U�����]�K�$�S��bCe��4E�����*󠣼f�|��;C��nH*o�~��x}X���p{o�%7%B��Ne�L��}rB{�6cǖ"G'���ZN&l�,:��թ�@�u�y#V�x��Y�M��4�:��,�D��!U�ɜ6⯍�j�E������������X�]a�Y���a��=áƷ�<�S����P�c)uc���᳻S)��Q����^.՜�����w��L���L��k?'B�!�p�9֕�)�W��B��mY��o���N�-zJC��=����RTj�F�k!8���r�͝�I�T�M�,��ѭD��8o(\��L>0|�$G\ $��8����vi��[ѥ�M�*�'�p{{e�Υ��i4;Aw�N��N�?����_�\��M�˳Ozg��J|��S�s�W�A��\�}rQ���M��dh�hn��B�*?)�~�O1:�xK�yh��6��~�J����;u�8b��p�E?��Ț!V �6�����#����Zy��5=d��K�ڒVw���^,���V�U@@��%�c���՗ȸ{�Vv��)J��5�~YLz�#�E,����3�X�P���~ʉ���Dw$�&�]��C�	�S�]QW��u8�w|^z�yHfO�7��7x����;�k��*�@VA8���0��!1w�[lA:��{yE�g'lorH�4�?%���+�/���|xkD�E�4��}��(x������{,�Y�1�2��Q�%�ql;�u�Rf����6�O�X3�`�s�`���ͨr��`�i�ؘ��%�G��v9'FM�{�����+���C*��^�������+���|�5�nV�^I�Q't@`b6o.�٠/�%��"�B�)��� 1�Q���yM��{�T�ZW��nL~�Y\��닧$�����E�a|�d0�zq�>䄜Bɹ�T�c2dt�=q'
�e�`o�)�̾���7�Ў�`�|�s�CT�@O*6�*Z�h�t#+�ſ������<��Ug��U)#`�_��� ������~Ʈc��i��!�?{�w�[6-��d8��R�J��pP�l$�%zX�6��VM�ԓk��:��gm~{�����>R�Vg+a!����J�Y�Qsł�OQ͞��]AmK�N����v���-�����b�� �r����B�@��%�"��8�G�G�,f8�ts?j���<�>.YCL�G��l.�U���j���Ɓl�W�]��f<�v]����z����m�`c�Qq�O`���_�?��r�ŰIqv����6n_Ӧ2�����'��&��W�|�:�ʨ��y�K�<Q��<�qm��̰�cza��d�w����r��\��=0K�~���9������D2����U�C*]���)��:/�Y%|�
IC�"c�'�!������^����3Sp*x'��)J�i�j���#[�GA�3��J���&M�p���v��Q|}�T � �p�S6
��%2�b.��h!/z7f�����0��a�_�Ea�6��J�ڞV�Zh�������w`yP��h��P
�hi�8�ٳc��@��b��u��b�S�*��\��;-��`<��݇�Cx�����j$f7㖳S���M���f@
EE<F\��N�f����2��<�]�
5�M�s�RE��\���K��{J�c���ф��/���x/����am\p�<�h?�?��y�nF�-C�ԱW	��Ėǯ�e�w��K�3����O	�Ԍ�
2WZ�
����%+�}zБ�=7� �okC%�4�\�i��o����b�ڕ��a`�� Yv8��[.=8�-�w�^ŷ�-�n�ۯ/>��~�!e��3[�A��b�SQ�}{l����\0K��  +�d���o�A���i�yV/./��������d��;wLci,�3�x"F��뚈�(ؑ�� ��~,��4�O��ţ,�O�3�3�+Q_�@������F�v�X���x�SN�����K&˟8B�a����:�����$�h-\�.���&�Vҙǉ:�/�~M*֘8Q�l�)��ܞm�Æ�|C0������ǢV³��$�9�`��B�]�ZZ�aw5-���Ю'N:H��*�ͧ2��sg�)�[�4>����Ep�w�g3�O}��ll�e�A�3HE\b ��V=��J�4[�m�M���ħ�Fb�Da�A�Ԡ�#\*��� ڻ�>A��]"j�NFE���ۘ�W�[4���p�m
�<�F�}*V�.�h��Zu��@W�%���*��{E�s���5_�}�q%G�s}�{�g�j~I�]�'�.>k��R�yV�7N*y{�1�e=����nȟ��H�ˡ`3 ��^��n� ���1���)�6F��O�g7�ެ.?N�d��`�qiC�T�u�x����h3շ|]�Jv� (���^w��ُ�h�Zr�'�y�z��u�b�:����%����w��EH��K�5g���X̻z���!Ck�3��gr�T�х�|�X0r��s��zʁ���n��c,=�j`�Q�U���S�â&�YfF9�3Oa;}Ih;����y�'&�[�Pz~�|1����!zMM�?���;������ںD�qǃ�������!F�^I5�Λ��_�j�%@��b9��J��r'�$�Z� ��Q:����E��<MR�����7��`"��g����>~�AYF�Z�`K��P��VF�Tݢ<ue�8��\�o
�/>��w��؄�O}��9��b'�iv9��#4�M��*���D�`��@�l���sL��__� ����7�9r4%.��z�r	;�KbJ�
�W�#�H[���+��u��r2�P��qe��h81P��k�
���S_�-s�)�`p��)�ۗ�%�e�x�w^���6  w(���hê6�1_�֜��Vs&K�Z����ĩ�K����*y*�n�Z�9��öB��5�������P5k��r��W��Y��:��GvܜJ����9��}�A�uGv���}t��7��l��{1���1�2<qxrh�TA�z�sE�/m̤>���Yv�_�7��6�����&�������	�8�O�kv����	������-�5�����e$=���� �Ѩ��]﫦g�~wu��9�7kY��p�B=�����2l$X�xȍ�8���f)d�^&qx����M�T7�
��q�^9��;���7�RZ�i�Iƫ��[���zԻ�[����.h�����k�w�;�?�B���5�GQځ�X�C�'F�.�k��+nn�ɣ��N q��JH��TmT{�8I�WۅCf��:�R0�V+�(_��Ѧ�D����g�����c��	W:Db�·P7�O�2�>4�$������]X(��y�B}|R=9���|����xv<��(��ܺ5t�j�X�*( �V-8���������N����]�oɗ>�K&6Kͣ+�3$�A���(�����7������?*}��m���]*�]>-�/��1t����J��N,���D<r��'����ɕ_[fR	ڟw\���|�3}{>B} ��䖒B�Oh
d��������y�1���񘞂��Q�i��yܛ�0�+[��vi�G��$y�9�MO��k��S@���������]�h�J����FH���D�l��:ˢݿ��dU��0*��;�2�,a��Y.T%>���q��b��6�2��#���\ِe���M�jM9���ڀ�Ш ��s'�B�����%�U_�W��1`��ǼH�xDYz�4�����E���;����Mj~��9꒤�fׂϮ�b��f� `��w��\�;.�N�����{P�(���\˪��BxeY�js���!a<G�-'� ���g�x�*�(��jbE��t'��b�#�2���(p���c��T�X��`-�Hbh����G]q�M��X(6�T4�m��?���$�1u�m���R���L�e��Aɮ6��W�2p��p�yY�f�Y�������z��f �M�-�@��j��;VD�YA��,��޸���5 <�$k���S�Y���e����o�0x��|��+Ji!���(�3�A7O>V%P�%x"%.��Ѕ�\R����O�G�6��Vw�׆�Έ\���r;��+t:�BE}��?����d�"��r��;����8�a�\�$c>*l�l1�{1Q.��3��Iֆ��8�Ā�w'4� ��&^>���$�G�^\��_ی*+�Q�d���@�aE��,���E�J�Ь������l5e�{>Q�8�k��Ӣ���N������'t���]������Xi��ArЩ&����3n9X�75�i��.�]Y��(`�����i4��?	�:���.��kS
m���oz[���N�:���+㸫��_R0������W�ܥS4S �|�x�����E�ZXq��)u���v*�j�a��I>�R�>K��E�:e|�>v�w0fO�:�;��[[�,�7��$�`6�}�#R�^ʤ�L|t���}�WYoN�	�ɵ��<�����e`"�q�e53HB���T�u�(A�!CB�;�i�i)�ſ�i�ۗ�}GV���&ev�B� [���(�b��_Z�r�������N]��޳�� +�Yڛ,J�ww�i��lK?@Y�* �v�-� ����qu���J��#%�ţ2�)��j�E���%c{��I�/@�e�o������$oT��Z7h�wT&D�2gAz�	a� �J�[���dJ�����*����j����M><�B�@.��jnt�\�0�m)*��Af�����@�H�Թ��7����f���N�,�-w%��B�=����EC]"�@}�(��k+����}�[a�Cl=�g�'c0/��n��q ߡs�N=D��q��(�@�	pbt�4:OxL'���i03�3?�I��d���	>R�!3�H�~X��/eJ#c�UT�S �P�`��!����SK%�ù��-S��ph�A��/ǿ�w��Y=_����	��ֵ�⸒S�x�����`ʻ����=�ż��@�3emDlE�;% �o���?��s�����&��b'�V�ءo���c�;􈫛Tq��L8�~��}�� U���4�&N��yt��"|uh�<GE����/>l'�������=F��,f:��;' �%!4>�e�EEA��X ����A���$M����U�k�g�]	ȫ)'�|iSy�X�mn|��XX�zʆ����O��Ã�C���s����X�s�U�@B���!������á�$���44��b<��km��<�^ϴ!�{
����ج����"��`�x+FFޓbk���$9��-&;|'�Q�t�ˍ��茐��e�(�>��H�����T�.�u����~���z}{����P�"�`��*��lx��%��[j¿Ƴ�8�:�
�V�Hx*+��JO;�Fs�4O�y�Ւ��d C���T7�����JL���]҇�^�6�"-��.��1�3�X~������U>�lY_3�a�0*3�>��R�h�	��;�i� ���a���3g�=��1�vv	[�<ZU��;>-4�bdjd@�i��B]�0��'���C��Ǽ%���5)vd~�(L�N\OF9�=��-Ф�<٬2 �4fغǧ<>�$�q!�ή0(�L/m%�Cw������
��6�>N^��(�6��+�!�ˆ��Dʹa��%�D�o�}]͖��!Ѓ��H�
X�mk��Q���^���ұx64�����+Ia�(~`�S�B��=��=Nj�},ۼ�g�{i���a	/8m�\ޯ=t8ʣ�eێ[I�ƹ�\`Ѽ����������`;KU/��&����'�V� i�+~�ߴG��1�i��y��y�u�4��3.j�
"�ۘ��F�h��Jd$��i�bpM��ų`�f��5������#3�M��_����c3�4��.�����Wz�Qv�д����̃3K�>��`?_a��brг�T#��Ijsf�
%?P0�?��d�$x���;y�V0�_d"�J/�<�K6.�T�"T�V8m�Kկ���sM�~b,m.t����.[�Pc����q��]Շy�| _0y�'=����`3���W� ���3�B���/��U��.���_�.��v�򒬡���;4ȝ��!����-\'��p��(�Ӽ�������td#���0��M3癩��U�l�߯�@�>����хF�����������c�	CHK�a��>�B<�`xQ(H������^��0��,~f�������f6��k�0��H?�%�P1У��}2VK�����w��O>�֫�����J�&Cc��K�<������t�.wmc�5���UN�=�Kߴ���ֺ
�W_�\���W������b�~GCl.�M3<Hh��<n�"M�á�a�&��{���	T����9e8��1Tp[ps3>�0�7��sk���bߘ�����o�^��e�G��l�I�����W��|"���E;L/R�6�7�-����$���I��b��-e��E'�w����/$�Es��sGxb�~^I��Zo�a�����o�I��O���a;#�-���,������t�+�k��JX657ys���=L,�p1�3Y�)h�Ddlo}f�_�]NO�*.I�ch �#�z��9}f�c�L=���*@����gLg�k�X?��S.x*y����o��w�Зg����V �w��l��˟1�L�Nf/���C�*��O;�3��?�Yy���HLz��I����~x����Ş���)h�E�a������SL�#�@w�|�ю_t��a����Մ�����@4y"��0UOt~���W`�s`"P ��>X�kj6�V�X�*��"��O�N=[{�U��%Z��}k���p��%�4@�m_{4|g��1��]���{1h���Q����]ړ���FG$�pH�Tz�;N�Bj)
Di7�_c�j�R�ߍ⨝�C~<o����v��;��1��@�a�Y�~<���K�d�����[�D���(�����駘�<%��\����Xg����~?�ç&��h3�z�V�M�N"o�hU7����	)���bx�3�E귫��۝�:ҳ�����c6�i�ۯ��Ғ��~�`d��-�-�H�'�I&��|;M�C�S'(V8)	�B�>����ǲ��c�w�����D��TK2�H�c�_?D>�}�԰�	��{	.�V\k��}ʯ���$1d��20-���e�0������K+��M����}��W�BTC[��|k�d��Ҟ�z1���� �|��H�Tl%7�Fo�$I��?�Ǥ9�v�[��}�K��ؕ���~s�����rM�d͙��/6J�%��秊��T,0�����\yP3��e�~.<��3�Ӓ��� �`�%�v�w�/� ʘ��{��?w�l�Ѣ�j�5�,^��m"�F�zR����0��L��8����n�(��IĀ3<���]~�c���H�媡�l�WUn?��{����9�5���h�9��?ڌ����{W^�,~F*B��2�_@���1���Ў�s^%�ʬf���l�X��#ֶ��n	�\5�ɉ�{_�#ҿF��U�LQ��߾�H r�4|��_dH��Īei�������H'����1�޳�(����	<E�4��9�&;�� J�-�C��L����U�8t�|>�ɦ�a�}��趈�U�	�u�|��k�ب���_��Jƅ �XJ�2��ɬ/����H�"W��1|�la*R��8�����m�AV>E���<�z�+��ү����{ٍ�*Q8W4��6 �yr�>۫�h���`#��:�Lҹ;��F�nz~��Q�q�؍�2�uE؅�I�G�*4��?�dW�V�ozx�ϭcOֽ�-%���J������U���?��L��pUSj�H��2���F���P�	�D���Ҕs%ʗ����Q�� G`���[}V7�'�R�s�<`F�,}P�{��'w/��Ց�|S-�.�f�̀�Z'��7̉��Y�:�>�:Ҝ3��0w�(SL���g��l�4̨���:���	C�k$���@���ˊ�)��j>a�����n����.�e�w�%��v-���!�ߙs�5�8!��@���X`FN����t[�
�-��2��2,�@�*"�lm�4,(�uT�!\u�!���E��*�{{Ƀ�ӝ���I��4	�v���[e?F���9�S׼܅֗�C�E#Q$��Rķ�[D!ug�JW;���n5|��'.C�:�ܘ�Hӈ�Ad{G�4�>=َ�pb6c���Fe��Ii3avTyǯ64kI-[��+.��	�ܯG���.҂!H�	� �5"?��u�r��S Ͼ
?�j��[>�?~�\���axEe�����@]
����2�U߷�w���:WJ*\��\�����Y��;�I�/"h��1�I�o���cv�D.��m*��رI�1��w�dZ���#cV	o=��L�32*�"��A� �����5�H�q�#�^���@�0�t��lJ��=���Vt="�m�u��Ͽ�J��H�mui��3- &�)e/�fZw)LhK�W��"��LP]ʴ�� :�k�^�D���:�H�k�@ɲqHW�	� �/G#%�֘��W~�rf�FbA��7�pf�"k'+we���%��<�מ�,!s�����At{����V�[�����}�̍��A@�*G,~^�>V���.k�PX]�o���V�Eϭ�RX�����i�n���<^h��)d�	�[~�{G�e4�=��J�q���%� e���e��×����"�e��Z�3�Be���Qi��U��4���k��?@p|�r콼|
�9���o�A�k�����ul~N�B��W���%�d?�=�З(��.˒XK*{�<J�F��9�_����7l�J�s >B<��)��L֝_�&�����y�13ʅ#�����߸E�q���H��NG�q&��f��⶯׼Ϡ"w �PcSG�!�c�Q�K#�ܳ�
��ȋ	3J�~6	��&M5�yW�2�a_�7�Fu��aQ�*s;ż��Ѹ!��6{~���o��p�˹cw�Վ.��L��jvM����ٴ(���|L����'��!���tp�ҚW��㛳��#Vp�5�;�cq�U�O�	��obg�2���X�5ZW�	�T�ׄ넊��h�#2,o�|V5d�V�d
ʹp卌M����D*�������f���9�'I:��ӣKm�Zԣ�d�d-_S�+�����2�JڅsH�����Ͼ3�����r�Z�%*��3A�.ܻ���9P��Y�2x�ҋ�ȎT~�J��1��w(ڄ R�Jt�uStT�4���U@�AҠ���I"��D9���p|%�͕�_�ó�0���Eۼc�*Y}\��T�r~�iLom�^ATܾ�:��'��1b|Gl��_>�����\�3���h�@�:K2)~^������ܥ&��D�)������;8��:��< 7�rh�!OJ�!i#����9�oGaY)�F���/�.�yR������b�;��e�&�⺄��'_�ל�t�w��Pn��l\��z�ظi��(S��f�����I�N*��fJ������L
੤�p1�!�I>��4�|�pl!L�����s:֕�s�Xv=� �ƚq�'5td��B*���O�q��`�=�����,HO
��=����'A��Sr
<�s/���h��Sy~�d&4�\&4��)�fX��˴��,�2�1�H�.��eE���~��l�|���kf��.`'P{�\�$E
��>v�
����*ޞ��ۢ�!�Zo�(�4�T��е,N���d��C�~?���=����S�������Bu���0�n*F���V[o"��)bI��a?),@ �oІ�J["'-Og�
��
�I�0/�GC��b��%_t{c�d	�>��� 8U�?R_��=�s����*v��~m]鬕e-����:��������`)�+���N�W��/�m��9aܛ���gC8h�ʷ^�~ѐO��~��ަ1� m|���6�� �r��� ����~Y�3�yג`��k�;�'���/�s���|�<gu���,\����4vR]�]}qd�����׆9X09��)Ζ)�=�Zy)��T�kf�Px��q��MѭW�����b�zk�S�]�0 �X�q�_�Ov���%�@��;�����Az�<��`s�NxVY���"cZ��SmߓT��	��2=��aiJ9�M��m�¡Ց�gowճ��g 8 ���&I@P��
��3���|����;�.��:�_�<ﶅ���؍M��4�l'����b�a�r�`h��ɘ�gTy"��h[�r��E��u֬�G+�ԵjBCɨ%s*03��&S��m�s+jX�co���#�
���N�Ꜥ��H��-G�����C��r��!=q�9�~��z�(w}��S�1�l���|Ր>�|���K��MH9��j���>U�B�wS��&|Ǳ63Jn�L� �Ɠ1�%I�MШ5����J��3���a�쎺�_e�#쯬fA�=>&zҕ?Q�Z~��"仜��<C���;��%750]���&� !�֘����(�J���4iN����n����}�M�?
�����X�NٽNF����3��jr��-��l�S�����ʎ�߿�2颺����=m-	VMQ��u�$�%��|B�d�9���*��}�b�Tv&7�X��By4j��$��]�`
��h�*�ڗ;�s�Uu�BYsI�
�@�;�%����gG.�QH�	����-\gXmh��I;2��i����4q��"U+�c��@v �(s����VN\��������?����TB\�:�a �a�z��N%ƳE���P�d<]NF���a�e6����|@;:�f#HMDt&x7��s<�h�|��8\��X:�l(�ۨ�0n�r���l�R���Ә�m`��U\>}Ë�>ǢY�)M:�L7$��oa`5V��u��|?�ՓX%�*F�h��l�yk|=��Dy�HY�E�cig��9g���a�{g��U����T����}M��(j߳���.�sG�Ժʲˇ�Ư�gZd��G�3q��HS�1{QNAaPp���=�Rݸ/ӁH�'̥$S�����8�O�`J�`�F�[Z��
6�Ū�>
fJ*��,pʆ<G��cH�i؛��~ba��R��j��3�Q��-�ʞ`��#���e��$5�����pF�Y�w!��̟�'�;�a����1�<�`j۩P�F-���ێ�+y픝+���Q�3��e��	�@ql����+��zTxz*�: �+���%��6�\��$�w;�a߳^��l%�$-�-��U��O9 &H����@�J����T��z4�-,Y���G���@�����!u�ˑ���E�5!����
�a[�����`�{~�����S���ïY*C�u�?"ņ���2�Z���.��x��G忞*�]_85�]")M�r�SLDA�k�H��ٷ�\,�׽��	�D�s�D%����JڼH���P������v�C�~_si�YKy�%��2�����4���ӳ-v��
�.@�L.@b!y�;��b��4���q�΂�0ɸ@�%�o:0v)�mCeӽX~�$�V=����(�h�Y��]~7e�qW��l�ל��"E�z���N�̮�o��s�\l�=�z+;�����^�~�Z.�š
уPÞ�T�_��@�QT\�2���I�L���O1Y�8*K���
��妔�Ǎg�9�c���P�mnV�]mj�t����װ�1I��y���߅p���҉����Ag�}��8��:2RC����]]5��D�R�KC\>��zD"O9�vNU
�������Q�A7x���j���_���^1��^����=گi6N�F����Vv�9!��6�Y3���IM-�+n����"o��H� ��.)�,pK���̞��(�vnSL�� T���uAӝ��+�h���R����| �1��\n��g���(}.���}��`���TK����m&�
>�����-6`��9kC�z��7���E���b��U\=kk���M�9Qde�eR�b|�ǯ�~��>%���J>01	țֹ����	ڥQ	�l}��c�>e�ud{I4Oly~�&�%#�d.+�no`T,��*��	N��/Oӹ����N�Cג�Ƙ)��������xSr�<V������Wq��ah|�����R�c �]w�HƬvld��s�t[���XХ�\�l{�;��������!!]��Vl{�ؽ��׈;MrhO;����e�D����\Қ	F69 c��sQ���ԧy�4e�1v(���WH��w�d)*HVJ�N.0�dW�ƅ|��Q�<���d�"�m���lQ�'ʧphY�^�(=��*���}2l������E�2��k��(��/W@�0�ձ�.ub��A�"=�"�ɭf5��cP��	��C2�=�W��D���6(����Z�Z��/X:h ��0��������
��kX����Ay0k�g�	K�L[��Ec�4�>�����3ٕ�%�a�m0I�m��i�d�W�)�������q�Y��Be�nHD�W"Mϝ�S����ba
�G�/������K�Nt
�A��Uv���Û�� 9����)���ֈp�i�'�,��������HR�
EA���
w�8�]c�%Ѡ��p� ���	�'����_1���&�бd*��Z�&|�rN@�%�([���qbj,���7�� E6W��qF�Ժ@�+E���Yڛ�~��_�/L�Y��2	T�~�/�*
f�������N���V��Ex:�ܣ��s�"�b�T�ϡ,c�"���S5����������iN}�t,j����s��x��%��VS't{?daQ,�i3f��<�sB�K��;Sa����꜔�[ς�����v�-�E�<B�f<���/M�T��j�����PW�\@K�SZ_֜T.Q��	'�Ģlg����R�g��bZyG��2���-VEױ<"~������j_�py�EQLW��B@XN�GZ[d��Wf˲H��}�.�?�Z19\�݈ч?����e�W�q�|�y�� �9<n�x��6��1kMhe�q^{�oDN6�^JcM��S!�R\/�{+`2��O����Z_��<�*䡃��߁��@�������?���+��Xn�4{���~9!\�DCQ����8����s� F��Yu��8��y&�\���"�~ k�<z��o�(0��S�;b�>��s-��NX3���Qߏ	jSl1U�I���^ȠJ'Y�F���5sdZ�Y�]��p������|�Z�)���e�$�f	uT�kV����rl߲+�g� �m�#�
��魱��,]
A-v;�]����Fs;)_�9��Ñ?ɰѭ+<Q��H�bD;��j�Հ��7�4=�k�\�����U�>um�8��k�|�/$�U<�ʙׄ���nx<G?��,�vD�@��10,�+ɳ(f��S��7����.͜�U�!�K��{ �ͅ�4��_��6�k�]��9a+���%�}�v���
����R
l. ��/�{Az7�LXd���.��;���q���[3����f�+۵�n���������ih���I�Ow9���u�z���p�k�kNSpv&�S��Uٮ*�9]B&�l��߆6���Ĭ�O��s�hn�#��[�������� �����:C^u:z#�<JU�}����c˨7�l�h3���,�<��Ǒ�^��zG=�Q��a(Q�B�^j��ٔ�U}̌�l��`7��ck[�40٪���p[���JG�jZc���Wu�0��aR��J+GD�\&��	�G�][=w����;���s�p��u�\���UD~ֻ��֋�`"nH�9Z-���� �X��v�X\^Ž$��σ,���Y�]�@O�&$O��1ͯH���ʧ���	1h^+�U����|�W{R�6Ĕu-C�,��9n�m�b	g�AU�eXX����l�D�f���u�y��_��)�1��ڼ��q���+cT/nT
oD��a��m5�Qf􂴃눽t5�2y�q�0�p`��e��\A{9bVioh�8��vB�laW�sjS��q2���_ț��9͍;/�f�#?-�Vg��G�C-xR�4�+�85��s�@ {8�݃iLF�X��z��>����T�(�5=`Q|�Q2n�`O������z��U7O� ��9!���D����@b�tm��w<��t��[r�D���K��:� �:gu�y@_�@��	x��ͱ�r�m��5�F�:�M�R;�G�Q�p�@��2��2|w7?��&%Ǖ�25X-h�w/H�C�;z����A� 8��U�g�)�묚��=��(/��B�M�d�[�d&�%7/I`���t�Z'��M;���� ���f�ŽU�i�9����'w�2T���b�9l������͛;s�=��O�K��E"h�pW�Î;k�\= i�q��S3��p0�!��a��2�o�ᡍ������dM����Zɬ=����b��xi�}ח�j.�4{;���:�@F��!Y�"�kI�����FG�u�^����hY`��%^��32�{R��k1�hVofhd���
��2n���p�=�?��g5�.����Y��梻�(3U�k��1k��/�h3$���~�FC1v��]$W�	7�����B5;V����O�֟�s�
��+T�Rwi����#�v�����>��@�E
�[2�k+��W���� k��9ʺ�#�ڎ���T��fI��=K���G	^C��5ȯ�v^��t� �S0�4}�?���}�O�	�e��/;Ĩf��5:��p�ek���¾M���k��?�.`S�y,�6�Lh���]�Q�|%��U�����n�8�1'&S��M��yU�s��J+b�0
�M8�q�����
���	���H�[�!Ha�-�����R�{CĢ�H^==�:mo�/���8���Ir;U1*̖��u����9��RZR��~��oAE��v-H�$1�P!s&S�H���mu>R��f��%�z�7�q����}ov�)�X��t��r{۟�bt���uY��?,򿶀8P�n@�yj2�k���6�A�ˆ��Gٚlq��FHEe1���I>�p(�%��>�8T��笖��u���T�X�=�����rUX*�絽��罠����TlzX��E���,�����C+�,99���> ���U��q������i�H�<����'b�����T��m�7G��@e��B:7��a9r���e���PM}���U8�S�kk����v�3���r1�0�3ʥu~7���**޶��D��G�7�5>U�~Ny_���Y5,��R�@;�7����7�v��3��s��L*Gu���������fP�&k����^?� "�����,CoPX)m*e��p$��Zo�[��nH�� �0d����D�)�P	�����M�l/:c8�1�y w�y�P��G&��S#t����E|k�X�)��� �ӛ$7Ξ�l?.�]�Q��&�_d֨l'�[底�w��?|m&Nb>'l�MU�=T!QJ�M��1ʑ�(��z&Tif��zQ���)�%�͔�ᐿ5� �:Ҹ[yRń������n���H�G!1i�'@�5�yO�ה4����y1ou�(�/?A�x.������jI�9"�;Dcm1 }`Ejd�RL�@���wB���оb�CuPz�31	{T�j�;��F[|����H�g�R����a�C�x�y�K=_�ߚ}�(��&h����������R��!ǐ��ʛ��6�J,��c��Z�v� ޴V�fm� ��M��v��62�����0Ġ|���[5��A�/^8C^���k�2Ye@�9S�t�C~��E�ݻ����b�o\{D������\?e�Im:���OK�<:�&ĘJ�oSZ|��#��u�[�;���*]�͗�=�[,�����˗���.����;=���[��Uc�Y��w�N�2��
eC��[�kN	'��&��K:�o_��f�5j����]�����Vs��Ag�K?5��=p&;��cwɶ8S��kR%&1�h���] ������[���r�ؑ�EQ)��-)���-�M��h�J�`뵔���hIz�c
e�{V�[����&�0!��} �T�k���
w��k1���TF"oX0���5����C��w���+���DM�_���
�����z��rX��l�
�0p���a%x��/�|���Ĕ��P��a Ɀ��X�N���&��IZ����[N1:���Z␑���Y�3�����̬��}:�ɴ2hNo�r�1f���}%���\<�b;IwJ�{#]'V�:i#6`%ПÃ�� �+��-�~7�y@���!��$�D��x�b���	�\_�4|Qb��ACD��H^�s�����)���Z�X�zѮ�a�\8W=u��dw~��(�O���Ɂ.����$����m\Rc,��EX/	�մ�Ӣ�/�.�r��zW�sx_u6�<{k?* �7��x������!,�էi��㝱ԧ.O�����"����+��ʘ����Ay��ƿ������>pf������e 3)b,�sy���M�fq��Q�5�AǒOHf�p���8�Q���X���i!�=$���0i�U���F�?�E�.'��G��X�M��\|23u�6�U���ZƗAݩ��&��E����vپ�e?����|�И�m��.��]�E��F�<�]'��A�9��q_�f������|a��̎::��V�:�z��2�Q(���@X�C��L3�F"�?�g.��>��lO/�r`��`af���w��<���v��%��P�ϭm���S�&���E̷���*x8��<���vj�\iu�ݦ{��a����ϸYRĮ�1�y�-K��3��n ��������4����=n��N=�5t�An@��9��9����^PB�j6Ҫ�y����0/'^�J�$��l��!:���[�mo�1��8&1hY0!@Ly!I��,Ub�bW��k��:�o�����t��>�u��"ı^�\8<@Mg౳�r�`Xz�[(�!k�q�{�s���'XP�x^vV�wS��I�L;Ý�F�*��	w���C����c!^1o��֦KwK�?�`��A|Re����r�mV�������t@�z92��m�*��܅�,���pQ����ڤ�alf���F��>�����-�ۮ�)�x�eƌ>���3��Rx�w�ᘌ�Ɋir����=f�l�z�Ǡ���
_�@��L1m��[�r�7��|�p�"n���du�[�eR�G���?�0LE ^5��Ġ�|�,��_��׉SL͹0t�|oP�~�˻�N�:� o?��5�lxd�/�i� ��><�ɂ�Q2�S�����yc���>j�%�۝���!jƉ������)�{J�X�d��6����nkD �4�}�/"~��E#�P^U��"g�I���, D6�~u�Y��m�;Ǉ��)�FQ���>�@�����jT��Wl�iT�H#�n?��n6�%z�1�՞�G@�qi+��k`�-�AX���� ���6dܠ��I�̴ �l����=Ē�5s����

d��Ѥ����f0�׬�6WH�bay	׽bi�&����ڒ��* si�$k�r ѹ�-�ն"L�D#�����2lw�AN��VnN��L
��B�N���k��YX_��ư0g���$QP��^9�7p�"k��r�����6�aX��MT&�i:�VW�M�,�iL��� ���,y���֞0^�nC�FI�h�{T��96��ѕ���O	%ɔx�H����x����D�Q �-&�0�ץ�.t>9�̋0�}~�vA�r��Ug�+��ᔰ�$_�7+R4��OVY7�1DO���o����IX�/H+Ai����Ϗ�8���+h�����}��%
ѷ�t���Ѷ`f����x�=�s3���qXh!l�zJ��'��4�N���.�/���	ɑ+B�����5�[�|������4כ|(���~S�j��sN�E��g�_Y%=5B~0H\�h�"�(戅˹������+�57� ��[X�*O�R�����P��#^�{OX�F�1>���r��U	��]�M+^�+1��������0&�YDg��A�
ƿ���6(�;&��v4X�-6*��)3g�|�jQQƬG`�u�����NS><����ISb�N�t��f9�~~���w��p	?�
�����[�7t����<6��4J3ƨ����/��	��-�_���w�b;[�Ae4���i�Xu�؈�n�$v����<$6��|/�hi�Ч�o��n:l��ܲQz���H٨s�)i܇�PA:E	������R���B�+_���� �>8���m��T;Z�j�Wͭ���w�9k`������!��]IV��q�@�d�q�s1���ʸ�ّ�_sk��QV�dJW�W�Rߠz���}���TIl�O�=�����c�j.�ī�=d�v�B�C��n����z"�+Ƶ�?-��N�.ޡ�]7O=�� �-��m����z��1��ZSϕ�OL�~�ӓxg�$�o�[6X]�	HFt�����]�̇��X���-��e"��ۀ䕣�܃�2d?�����? ��e��߅�/�E�y��v*�6�.�쒟Si�*�a�@����^wc��5�T�$^��������:�+�z�ˍ��`]���t��z����紨�9��=�����x-�_�`f�䶌��zO�����0����Ʉ�ѽ`R_~����A�V1m�>�{r�⒯"�z��VL*a#��w���?�G?�Crv@�G�h�t*Hi�pK�!9�熣٦���.%d�#���f#9lH�Z�c��^̋�*�R\��b�T��_YUJ���~����	�U�a�킾u'�
G���whVJ���ΖlȨ}����cI�>v�h�볞nm>��D#�*����@���]����GԐϖ���O�3g�"��Rǝu�Z*�jl1<���0�δ���^��xj�����nM���R�kX9,_w�Q����	�B(�)�2X�v35�S6F�6���NI�/'\- =��-��Td8��-O:�D�T)���Q�WI����D��r���839�����@���=��}!�\��+�����O7A��	l��Ӿ$�����;}�#���Vio���l�tx�����3*&?� S҃4?)�	ܮ�q'R�b�V>^t�!@�'�U�{��B�����@2g"� ��H_�_�\g�IS�ȵջ�5F�TC��8��j͢P'RMM�Dr�W���zȹ2=�3k/���Y�!l��O^q�6�)�C����>�/�-����nL`� �o�bm�31U��L۩9v��
m:�����d��M0��()��^�_����$��͗aH��� M�0�� /4:��n��!��}�%�!A��S�L�U
��yUi��A��L1��B�«ha�z\#{������#���z ���w�a����ul�p��w,͎r,.k!r�}�����`!�+��+���L�l���l��j6ȽO��Az!D�=��y
��'��5��x�N'B�م��˭����Er�N}g��K�`;v�M5����4�����TNwa���&c?kɻ��y��
�'�5�ֽ~g�.�z���=��(L���X��3F��R�cl��>��S���x5�I�>��b���a* �sX�#wh^ � %ʷ#�/7�2���?�Z�ZC�}E��I��~�b���������1�����4LR��[`6BR��11�CȰ�/��h3�q5oG(�8�$��`��vX���I����D�᜻posʷk�(-���1�P|��^-���M�f��3�*9�v�/�=Ĩ�\?x	Iy,6�C�~�)6B��-�W2MQ�s߭+��=!C0U�
������G�,a>�K��~�IW <T�_�����(>������i<,:����8�a��+w~U9�1���~7�B\���[��D6#�+� ��7�o�p�tǲ�Wm���twT*��[-�iC���W0���# ��m����67"{���#*�CO�O4w �3l��C5�>nĝ@��tc�]��襧�:V�y���$����z�7#�MW��4��q�{�B�Wg��6���'hAx{�=X��>?ts�	b~b��S�=� A�R7Dr�"���o�(��Q|)4�<�����V*��
ii���0���!ok�����,BH3������*�g7U�[�eo%xtz�ǫa=W��/�A�R�� �M���f�ݘ�����?]�X"O��i�@Wy��'����a'��+�qco-�Or����w�g	��}��M V	x�TI�$-n�����%s;[p+�gA�F�b`D�9��vw���|ÿ� ����ILj����L��:��aQ� �'yP�љ�Nz���,8�.�V����<!��Oh��l��@�֢y�g��3ڭ����@�m���>�U��6��<lvO�]u��T^	C@9�u7���? �q�q��R�b�˛Kȴ��*�}ð�����#'���P�	��x�X�YZ�g�����m�<�46'P�r�f�J�?�o��;  P��p��X�,a����MM��Fr��'.s�W}϶���<i�J���-��(�x����4j�����x®/�J�cҞ��[-�]���db�p8<��y��@L���Z�M��M�ю�QV�C\���$�=�[��8<F.�����e1� �'����Z�l��Fbe�t$غ&��εQ	��5V�鮥D3�x[B��ζ��6M!�mOSN�މ C��_�)c��l���ژ���_�t,OM���1��(�r1'tq��l�w��`�_�#��t>�	w/�2��EWt�zN��O����� H6�ڬ)��U��˂0qu�;}�/�Q��{��-gKb������֋_HA�g΄��gi�Ac"wUB��}Q< �}A; AB	Q���J���|n��n$�~�j���&5�n2=ؙ$Q|����H�=���S6�Ln�<$�	ը�2�WsȆ�n�j�|�W���9i/�����{%��A�-�T�;'�ȝ��/�\�����s�]�*�Z�"T�jÙ�f�sn�Մ����1{�H���ݔ�f�r;��:��r��]g!��>C���b���e4*�o��P�r
i �QǀEe�����2Sf@Gcډ<�%G�c���Ujg���>M��t$c�bT���GF���`���
c�rC�`$ɫ2�͠�u�O�ϞWl�D*�t�`��uB��#�A��9�s��>��w���Z�j��mw� ��� Ea*I0V͉��@�Ĭ�3� ��7��P�>d�����9��9	���*�Q{ɭF��e|�=�&3R�i?�u��S�z�{D{7!<0R�օ�5�[8�.�H���p,�iڢ7�B����=O����g�T�\�d^;�����ƯE��V��r���2��G((dN�YCDh���(�\�߾��ѣU�9w����,Qٯ�������L+������PS!i<�>WRz��jQU�l~�����Y���&��L�z�m��.���C��"���N�2w.�f���mҥ��t�}���ݓ���=�lVT���3 1�����Z�w���O\� ����ٕezz3��m.�/�7�?U�O�.�d� vI�K�3n*��!C�L��0�wYs�ؖή����
����~9E�Gm�������r��W5	s�?W�i�Wr�4isWe<��y�+ܑM@g1gUzI��w�Ho�ȼ|��P5peyvz딷����(��%�K�]e��0�פq�	��P���&������0�/D�E��۳m�>7����U2v�v߾�d����=8	����̳j�-'8����)"��rLp�Y.0����qyDՒnU`��7��}�*��dl���6=v�(G���]붽�w~��O,_=����r����h��`R��A�oH�ӠG����߂0=���΢y5���7(F�D?�m�U�o:�D���|��qo���l���#p���;u+�r������x1h[���{�F�^Ī:Y�V�0�0��C���Ze�t�ur�SG���K�$�<Gթ� �k�ّ�	�f�?N��������<Y�Z��	l
U��\u�(E� F�D\(l&I~*�?���aذ��%���)��]��D��V n.��.��

 6�7�Ɲ�%!�H<����N4�����s�PYb�X��#�3`��;��7��J^��Cu(�g��5�sz-���C��_NTS�M�����Os�͎��u��./�㽋`��w�s����'�boO�
k�#�D����w��{^�π�#��.����n��M�F\�(1>F�_ޚB��@�,h�B��{�0�(\D�Ո�9?�;������������t$�ú��zyw�2,9�l���EР~�o37Z�,���'iJ>/f�y���\ˎ�+JZ��3��7ޙRo�sBA~Il���=�2E��H��I��f��k�'=a䖋�°�9��K[�8>w~U��|0���mq$��b_��ל�L�٫8�Eh�K7�ϝ&�>wa��u���e�{����L��~��e���\=���#p�d�΍�x=�>2$L�h����)�����b��h���7c �����"�FVV/���q���q4�s/���@�A�c�T�VƲ6�;J�b��*0�����:pQf&VS�v;Nh��e��$���y����q�~Y�H�Hm[��z����H��8NDH5M�Z�6�R����-U'�]��ԧyX�a+���Lz��o����~ "6fr���"���\z��/ճ �?e!iT<��^2=�hS�@%~;CB��3D˝r�s�r�dơy�T��WldC�Z>�ͳ��S�8����m4�>�fq�ϛsTc�֌TE����>;�P��$���إ�3J���7[�N�zw>�)�$����"��m���L�t[I��f@(h2��5�y&�Г�B��Ao��V��]E��ʌ�ʴʤ��n�f�ؾ��&1���q�l���'�Vj��cv��)D�c���X�_^��݄�w�M�Wk�)(��a�F&E>
�J��hE��c�̿C�n�t�lW2���W�����t()xWx
���X0�������" G��G����i+�R�V�ف)�e�6����.������I�� 
�*=��2I���H��U�5*8�`K�l�雌z�� �NU2g���Z!)<6`���u_?f��"A�Va2�u/�H���@e�^�	���4�=_��<�!�^�����T���@׿��1*i����#�p&�5H�b/E�J�#�F�/?��ĝ����,��C��ۼzŅm�V� E�_56Xw��l�D��t�N�������_��ܩt{�D�V���-�wj�ct%�t�H$�3䜚�ջ�N�%P���7ů [��xG��
�h<yQq@8����0~q��=]�k3	���ߜ��I�����6B��H#�<6�S�f�����5ǭk�G]���9c?��<�=&q~�m��T��1��M�#���-���P�2���=}���}�,��}׳Y�<�C�~���W��\p�7�f�����`�yS�C��Á��p�T�P'�-��젼�5�k�N�ZԂ!Q@�?ye�MMw7��&I+`y� �߈9����]N��Q[Y���m�A��cw���{���E���/M=S��j��N��L�p��[�9�\��Y��w���$��`C(&�nU��B��t�Y��WL���W�l��k/�ti:����=�"���;3�51����0n8DC!_�m#�\C�!�9�,=�'��\ٌʌ�������>���#t�xDD8냫=%h����r��݊��	����i�����O�+��8�s�� ���{���]c#0.���<�c��,goO�>�|LT,D��2:H��E+.W��2fqyJ����&�Pԛ���t���Z�Zݐ~��f�Vz�S��P�k�J�QYS��.'�s����[�略�ǆx�H�aVg�������y�u��,����,�)���f�
�h1�ZeS/la�ˑ�k��y���'�9XưU�6ʲ��XO�5.�= �P~��o�]9��-Л�|�c�-�5\96��2�=UZ1��L���U[���H��r����`1�	��j]vr,���C��\�?AbF�[N� ��`lB%�:J�X��(����&��]LZu�YT&`�p���N�D�p;���#i�.��ܭPO�Pi���5,�UT�%ʇF���U�J�$b+��<?�$�'�ƚ�N7�Xơ��'Lؠ^n�1�ܥ��%�(R<����R��7��x��Ȥl<������ED61f��0����6�����~O44@��(���gT�аG���r��-[P�u2ъ7���&��S�-S{[����Y��w|N�g^����2j-[�9��U}��VJ����]�M"W .�4d�ꊘ�~�a|���o�!´���8��o��%"҂���CF�߽x�d�A}F��IBR―��]ox:�+T�+���O�1�񡨣�yB@��m���8'(:�}��)1�K��~���=9����z7��٥��ڝ���i���́��l��!�rb��(�k+�ӿ-n�;H��	���z�K�3�)�/S<IRA���|�g�q�z���	
���s.�+�#N���Kn� �H�횯E~�Ȭ��7�em�n��^�ʤ�6\����q�:�0�� ��G�HD|�6KN���nx�7����H!��B<�D��6����_@�R���|������֩oY?��6)R&�a��Y���McQ����/�Gσ&��1��//����с�mJM6�n%�e|�Mr��e·��n�cr����Ƭ3r"zҚI�*��'�tr�4�"�`���B��k�IW�(q�	�1$?Ck �G�%?� ����j�'0�4�}����6��-�G�9�����lB��M�6^�*C�]�8؎J~�\oJ�/��M<�b|ؔ<;iB�eU"�
�u+����в8pn<�Ӆ��b��^�ݪm��e^�RJP��[�Qc�]O���n<����:ֱ���ӑ����v4�4M�X�i7bʠ7�~ ,�t��2o&�KXjsj��o����-�c�����2�d$F��?�3'�a���nCՖ5g�O���`M��S�D�3!֎D	M �ȵ�tW(���G��_���US��\)1}ҥ���eAbiC��ޫ�q�O�c�t����Ɠ�O��W�`�҅{�<bD}Rg��#�q<�P[sȿ�
�^�&�n}�E������\��<�lZ�-���G��	�+�J���q���=4�})�(K2+�G�^Ѭ���������;����1��!�܋�ɉwf���"DN�xu>AY��66�[�]�]p��QC;=A^�丩�nm߷3G6�i�M
�$�3q�S"�'���:�f�sgv�̈́��������f0�ˊp�z�US�Ao���6�+����u���o� �d������5�f>���q��5��aռ���J�i�A/��ʕ�d����:�/q����r��1C��V��}�d�;NN��[��+���Ux̰п�^�u˧yuN�D��{��Ҫ$�4B�Cb~@\Yd�dT^W]}�;����6����p���ǆC7�VY���Z�����G�W�0��g�����%�_���Z��t���7�ؘb���-4*?���h����D��������mC�7�o��I�F�źF|^�� 9����LYx	�L|��!Qڄ�']��3�Ks�Z@3MO��7�,'��jA_6���$�y��W�[?Z��R*�
�B{����B��U��7�iśԕ@�N00A���V%��g]Sz��U�c]���ԑ>�s8g�ǧ��IP���}��iAm����;i�B�g�U���L�S���U�����5�C>J@ڈ̐%��찞�<���A2�� ׅY�����>Q
s0������[�<����u(���I�?СN�CjR N�ܾ0��>���'߱h���ؘ�;��5rد5^en�V�0VUp���9���3�~S3����]�*I�D�l�i������C��h�+�	�T>,����[ڎ�vr�/�\��g��?�+�yb��1�VCN&>M�¨�k�%��uI;t��z�R����nS�g�����4W����z(���R���� l�m��ʉ����(t�b�E-�&4"G�P��}]��F��*�)� "b�L����e�r��7�3)�[�τV'�*'��h-;�
=�޲��:!*���¢��S�PJb��-+���)���!n��,O��8S���k͎V�?Q�������b�Ή�U1�c5�}�U�Uv��g?�c��OA4\���)�(jEl��HP
��6��� /��QD5]z:7Ζ�P/� �Lv�:Z47(}Z��	LC�?m�6�5�V�j��I��rN%�0z�xt����������M�Cq�Vx�/��q�2C�7�yZe@��9� vU�S�R'�	]�x��;�(�P�\8*�ֳ��0.)}di���6"t8���V �@ ����Z�es�u£.�<ΛO�B�r$��ȶ��+����q��N��ZZ�&�F��#/3N�����<�R�������S/}R�+�v�.ӳ�K|����M�	A{/�"��ح���|��)�����S���]�֡�9����R��ZA�7)����e}P����#.��K�0��>ч���.�u�x7Q��U�K���v��o��Lb��"�b��U%_���O$M��7S��;/o��F���r�	��m�W�-�����Z�̬��@Khr ����� ��Y����ӽ具��8=ZA_2#�RK�μn��>�pvļP��D=��Mk���#�ZE���<QaO�D�e�K�޳�s/���9y�4��ޡt�s�f� (���d���wś���H��οɺ<����_�x�rD���lx��	I��k�纺�2$��Y�8+VN���Y'C"EWvM��q�a�a��X2֫հoFR��}5�bux��m�)u�H�`~�0qR	�������pF��S�(�EkM����8������AW��@���w��p�n#u�����Lp����g��IBxb%� <P����� n��_'�����~���ذ��(^��j�[ ]oI�9��35��� q���^�RdfGu7�����c��< ��d����!�Ks�O�c�K,>�an����$n�Ϋ���Ec���/��}|1}���@.rI!�9�w��H];�M�V߂@�1�z�g�G�9�)1&��Do-`
�k+����y! �:�9��']����ό8Ey*6����% ��B�s����Mw�a)�c2�����q�F�U{�&�����*8J��3�����N�� <�p�[|2�P�d��Բ�K������4�4�g�D9iDK�ڗ�v�e�2�����_Y� 9�l�{>� j����*$f��(�Џ�y;1�p���C�`
K����s���u/����Z��3{&���YU`ꏬb���Ԏ�'Е�H�M���w�_3ഽ�]L{��ڔ���e ������4�x◪�{���!�#�MO�̝� @�9���Lә϶��J�� ݓ��_2K�6�*��i�{?����q�A��=��5b��/9�Q[�Q�ym(��������@*�Ǭ�-68'��-��	�n���=���U$=iBf��n�1��zD݃�o�N��*����sZIw�U�n.^O�Q��z�]�%���T`5�߂�B��+����h:f�N��x%�ɿoV��r�k���OH�t�,�qQ��_�%��C 7�	#�Q�E�z�m>�"���Zg�OOc�ʅ2���5�!ή�Q�4�;�x�	�U�f��N�g��ׯ�Ծ&q3���X:�@�[���`;�By=�׸m���@����I��"I[��wSI����F�8F0!��\�*��j���fmZ3C�v��GUj`��*�*�I��b�߈��"�U	�_�ͺĘ�ܴK1j�2E�Z�nׯ������-�����-,�h��eyH��5b��7wY�T�Y���+/K�P���T����;n �=��f�y7±J��Ih4���{�����$Y<4��u}ffou���g�l��{� ON�{S�P��D5{!��t��&
v�@���u�\<�Mbp��b׳d`Y�e�{��z&d(�j���"ʪ0�E_��"������-F㠖5�c����9!V1&'�{�x������=$�'/�~���,E����
H0GBnc��DoO���}QS�"m�i<aS9R����ciG9����>�0��If�F��4���Ա9�U��b��H��۷Fྀ�����}�`�yʵ8$�o����,o�uA�gk��ר\0l�#yq,";����_��,�p��l��_�ڙ�w��ƫ��]��c~_��R?�b@mٳL9;�O�TW2�߀��]�T�ܾ\"ou-9$�G��PE>�;hd�	~����PsZ`h�~Cm�K��t{�G<i��ig>5�&�^2�u��9ý��C~��8y���~��'|�k��gڭx��� �j�7A�:�sȊ_ϛ%/��M{l���m:�ͤ�r���{���R�h��
�1��&P��.���8�3rˡ��qhI�W���{����X�Ǘ�b�~�,N�-^G3�I��پ�J��n}�+�ٕ��$��ح8'�@����oN|�e���E�F��b�EzY�g$ ��	�Hҫ�b �к�L�@�q�{"J�"��9����xO���5�>}�`N$��3"ʮ/��^>�εgF�>E��a=�7�'���)�w4x���j���._{�R���,F5_���u��=���T���N�SDo����7u)��q��|�n�`�61c�~�܊/��z��;�]��������4-��Q|�}�I�S�%� s��)�� ~]�C�Q|tW�g�[(:V.�M�r➍J`�+�0ҧג=�;n
�������b��x��=k{;�70�c���m\)[T����ւL�n;E~���fu���w�\�[R�=#���J�xa�q�.G��X�3�����t�}�S�+1]o}�}�N3�4�`�z��vDJ���)�:c&2�
�P]��5r�D_K�Ђ�u�F���^d��	�Wa���t>8R�;L9��7+U	\9����3i<�ٴysT��9�&m���U�&���%��Ԛ�����5��ٻI�VY�d6��z�?�Je����"��ج�
���;��������<z�M���Pٞ�аF~gE.vM��<�g{�@���0�Mm�Ϋ#��긙7���`J!J�ЯMA�!�fC��+���4���� �A7)��F��� 3	��̋]A7�w������1�Y���M�K-�r	D���W���U�U�j����z����g����|԰�'0���Ч}��jM���F���<���Qs��ǽCP�5b�1�d�Q�~Y? ,�bL�.�9�b����Ֆ%:��&�^|S�"���?H�>�xoW-U��˟Zu�'({�焃��#�ߗ�I�4��RR��i��ƍ?@5�3�O}�;��Ю�&�b��M���L�sE��Yc�6�]ʉt�e�':������&�ÿ|��]h�k�.�R<ONT�%̓�%���g*�U��ѣ0I��R����N^7.&U�>7�5��+���:T���I�䄻�}����cgց�i�%V�[z�`EI�uF�}�-�Mɟ�"�3��7�j-�o�2yߛ��J��
�!�E&}��ؗ�p�u����Q�Ѵ����@Un!��ۧnܚu�/B�4s@(������o�;j�l�6���`�2��ԋ]�ҭ���#��a�Ji�Q�a��lFf���p��痫,��5f(�؝��m�$r�CBka�|K�R���v��Al�V��|0Yp�j�ۣ,1(��?�x/�����uK3�Ū,��6����t��|�z��	96L���(r�|v�2�_}q���I`�rt�Z�:��%[�2Ǔ�pX�S3"���r4�DL`��;���v��6-�؂�B!�t�w~�˻s��r����$ƕ�R%/E�jdD��䉼|�kY�� ���I����]$rp/�kt��_2k���u߄(ha~4��'	��{/��;�.;��-V��}лJ}���*�;X��k��7�J5�F����y�lB��� ��� �p&��tl�/iX�U����7��[���}C�IE:ᑙm�胭u�P��>��hg;�952>�ςZ��w��w���C�L���)��(�^+T�F0��f�.��4���#<4��
�S9B��}���R�TD�q3ld�!�4���1�ˮE�1�r�e~���l.�(q�N�a,�j��ؖ�/x��s���%�l�D����o��dB��O��ا~F_�Ra����v�A�}U�hs*4hs9�p��:<�|]vĨ*������n-,�(�L��׬9YY���Df�S�E"Kgn�C�v ��r�\��@�����_�'F,M}Ӡ)�����ҁ��w�|�6|	3�)T�E
Dc��+ZK9�Q��a��`¬7�t����\��� ��kr�ه��r���y����ٹ�SR����E��e��:(SW9�PK�>�O�γ���[����e)�?"���IO�Γ��@D��8�0#;�����7�wx��WWu�fL��K.K�-�1��l�p=���<�{L?����H3<%���Y�i�O�JހRO���-�qx�JI�.!a��+�j�����)��Js�P�)�O�fEH�ϻJJ����6_(2��=VdS�������2z����%�;=�8Ue�Ϝ��ڡ����n/�8R��щ.1f�V�L���|h�r^�ok��̃2pd70Y}8ld5���Kܭ�ff
qw刘m�����H']l�%8˒+p|���c��έ/g;����h�gqN1q[n��e
o�ٌJ�+�/lX�6bF��j�b�:/k�SW�3�rH�(B�Q���!g._涊���V6e;m��\�}$�-�5D�7�6:�0��yg6�$I-n�I$n�f�r��Y���4}�j�A�-����ڠ��mYC��O�ٹN���$X��[�q��e.��>u�d}���0��b����D�fƤQ+`eeI���A��O6�)�l��m\Gp��BW���c��������TaR����@��z-��XJ�����Y�_��;�	4���X?���2ձ:Ё=Θf)�j�R���ĳ�I;R@����+ey��UJ��;[Fhi�e�$t�R��' ��4b��OM��/%�@����o+Z�#}��
(�(z���u��d�Ra"�r��hZg$�J�D ="^�.���݊����Mª��(+7=Z��Sw�6`$(s�����p_(�dΊ��@�L���*8?@b]d@����_|�I�[�P��Ǚ��Wf4��U:X�A��)���>����������e��-�,J^P"�fC0$�⫍ _��^p��-�����&�.�!"wv��|cM�l����
ݨ����̓p���שּ��ƺ:�y2�h?��S6�:�W������U���:���%"�G��SՀGc_��.����[5��� �B�3x���Î�L~��=8��=�-L���8��?�rσ��1�.��j���ᆱf��l���t*�d`uG4����n$Z��%�Ƅ�Uat9��H�k<=y30��M+�P���'���g�����W	��oЎ�z�� s	h=�d��/]�G�M�g��<�i(Ӵ���3�a�{za[|!	lVDqM)����<���2���P��P,��_!UG3c��z�_�~��<9��i����[E������}IG�/�΅Y3�����`�sq���4##�LsU���p�x?<^�L�p��/`�L���{��R����Am]R��A��M_m%�|:��jp]`����r�!���i�m�/�l/q1�rm��$F%o�9O����o�\��2�o��yf���>��B�P������� �fY)w:Nu[3�V���&ѮM)���}���F�&�>}��R|�������<��л��LD��� �M�FǴ��|�7��W��P��V,vEȕ!��x��v���/�����. HM��W��uJ[\��
���A�4:v�3��n�ʘ�񎼋�a)�}��!�"I\���6�`���ߌ3������%����J�R�!>��Qԫ5V�0�HY�����֛����{������8��=�4���W��j����FF_���p4��"��c��UY��sE��=�v*2p��?q�����/����[}�X ��>�=W���DmE��T]�Qw<tr�?��S��Y��٣�FA�(�%�[u�`e�i%3��78���9�9���{茷b�eh�Z��6Pq���#���x���g�<=���������1��}�m�c��� ,�����Hn������r�`�?���,�j1�S�P�{��Q	�(ܣ@ /S��D��'�1�7�HԘ�r�5�[��_r`�����u>�0F�1'�8B3�����5�(�����p��G����V7奞��\\��'EL�'��,vם�
'�����Mrʨ��9��F�r\aF@��47��$i{$Z���i@&�4a�U�O��'Zs���4I<e���WySǯʼ�x.rb������uf�I�*x�'샜�!§�v"���������W��#@�M�>��f����w��ҩ�Yև౺m]Gp�\C�8ۍ
�
d��|/�z��Dc\,/�"|Lry��F.mP'A�)�����Ϻ������P��ϞF
I�W�Ç,��X�~��zؒ�1̮�y{ʷ��3!��V>S���pZ>��S�
H�!��t��/�'4v]�q�f}��:���8�t���Y���o�<�S74PXU��m�c�d�!*9��8o0 #-��m�bvI�
(U8�gj��_!K�"no��"������Z�!�C�7E�V��aa����/�^Vؙ�[��b���4Y��`Fs�fU����2��*	��^�D-��]��eP���':`w���*�J&̡���l?>K1�H�%�<.�|��1`G^Y��ҥ�4�-��X����?z��7.�PS���ɢ���	���{� ��v>��Qk�י��}�K�a�D�Y�[_oG�̫�V�`D������,�4%{���S�rD�4z�e��j��[:�B;���>&k5�j;�$I8���JEPaSd
G!^�,l1��D|{��!Å�A�;����"80l�O��?�cD������!���Q<+}��IRO����ns�zjn�g�_6K�m�{ˉ����㥊���ޭp�Ԙ�����$���U(�S}*o��1
�Q��ճ������:��IÉ�K���`��;�1x�;��ʴZ-�6�V���Z�d�����<H��_���!\$� @���ێ�T��D�6��M%^�֞1��p���^�u���W����ۦ��t��r���E
x7~y�	���Nn������%�ž���}��@߆3u)�$�@�ݢ����e9�;���mg�*[�1��{��0�Wp��,��P��	��"�M̔���>Lk$m��e�|-\�<5���H�MJ���B��&t��QH5��|�q�ZG@�x��-��>T6�R6kb�`�:$F�sѬz�#3��$t�,�oĖ5ߝ�$&�rX#h?�/�<��*�u-�N������I�]z��F!.E_�5L������_�w��n�+-V��2���k �"hI���]�_*=���^��j�,�yI��xD`N�]aA���]A�Su�2��Q5"�]�l�6���wm ;�=�M~|/�(���'b�CO��;��FՉ\;"�\�R�)�bN��)�?�������Y����I�
���E�O֌���@����T�g:Ms\U!�,;e8�ORޥ�������}��
���-K�0v��CݮG0ʹ��e��ͼ�C�LRkj�G�~��"�5�$�� s�G	v!J|�˗�R�I��Uў����]���*gN]��<=Q�H�tEvB�u	H��`e��`u-
��t��5ց�����jx���#��"�e%"I1}�dW��L^� �6-.�ɏ�U(��^��M��7�d��ń�
ȣY��!f�r��>B�Nj��1� qD��2�����?���8�#�g`�Y2:�W.���Χn��[�6֚�u0��F��gl�K����Rw>�s�+E'��_�*�F���c
n>S�w�E�q/���{>��I�p�N@.�L).h ��hb�(�����5��H'�3x�O��U�1U�$�t�3��?���qgJ�oKG\�o�vf�ි,+���F��J��"��]o:�-��?`�/! bo/�J��\�r�Ʊ<�m��6ly�A'��A�V�e�M��Z�0a�K?RK�t�W��3u�iOb�h\ڷ�/��gӳ(%7����BHo
o����g�E�v��Ճv�r7\ ���C����r�$=B��)a��G�h'��+�a�-
�������ބ:�����H�\��^=i��ABB{���ڇ�N�=��ܯ�7T�O��?.v�g�����L���8nc��@[���m�4Ǻ-$�F���c����{Nk�~^V	.��#1췛
�"�%����XS��
�U̹����:B�:7�X��I 3^�V�$�Ff�|@�Pl�4������b(L�=�.� '���F�1�@~��d���͒,����+��j�_�"�3zB�a&50�M��\\� 4�p*�(��A�R2飲�1�x���0��[_.��(���j�9����-�e�?�����X�O�~���z��[,�*�Z��L���<�ξ�@9r�(��`�G�˨M���InÂ�D�Jv�y�1GA��@8_B�'��ﰭ�{R��*��:�-��	jk�8��F��,o�'�L��r����B�3��N����u�n��5~jz�B+���p��� �(��%��$9s�濳r��J���D?Z�9��q��bO��1ZF �~df���׶讱8}��o"Φەd����fyp��^��@����d��~��:�i�A�4e=����i�S���`�+ � ���HZ�Fb,�����0ƽ���x��>����S��D��a<�y�=��&�C���k�	K���O���������Xu����QJ�{u�,2�`Cr���]��AzO�'ǁ�5<�=7�e���-����d�Ȼ�Q������@2J�g�2�#�����������4l�Qz��6�=�7������,8?�GbP�VtUXG}ƺϚ����h.r�n-��#���2�2���hQ�+,�D!�}�$
=	EUn���?V�[��,���-��ѱv��5]{�<��Q���XƀG�E�iY��[�3B�ݨ���t�֑�P��<���F.'��n��ã)�W�ri���-
pZk�ˣWƺNS�:T��{�\	���8-����f}�n��Fߩ����*韹�W=��Ic��=e��ʋ�I2����%�[Mp@_�Z�n�.��s����S&289�V��kz�A�T���Gk�p[5G`���=�]
7��b8�WӰ�;�Q��ɟ��Rl�=�-�-��{��K���O���g����X���^��n�A����iN�)���iK�FRE�e)SN	��������u�U�v����꬝�j��m8o�S�O���d\�nm#�F�Pԧ(��d4X��+�	��	E(�!�>>o���x���RA��d�X��U3���&;C�CB�5B+^.��3~�X'���@�J�	� �=�mqW����t_7Z�����{O~�U��E����;�P�Ժ��mu��^D�v)}j�Õ;v�^�u�������G&�����ƿU� ~��j$��؅�:�#4�-���c6�ϡ]�@��"	[�|�ҧ���%h����������m1�F.�zo�
Cz�+hQ�җ}�^�0�o�9*>u���D��\-u��q��^h�������2����ٺ��D��F-Lr��ʲ�^�<�r���=+��؃ܘѷAq6�3�J��vC��)�I ���@(�*lmb~C�<��<O3⊁�j�*�nq��:��OO[�qm�o3���a��& �P]��Nxɝ&�
S����1��?TT��.#�|���ۯ�:&�c���c�k�jM'w%p&'C����g��/��*�+��30_hdM��ghv���~G�-!����-�����̀���L��I��ld��
m�$���]Kp;������#�Q!�4I4ۆX�\�?x���~��,�M�i�V����Z�ૄ&^��ˤ�d)L��}�R\kɕ�||�� �8z.}
�aG>�Uc��o>I_�0�K��bL9��-�[d9�Y�OԊLnfE�{w���"z����J:��,��3�:HZ!!�L��g���0.c��hoF�2�E#I���Ո��{y�!��n��.��fR�aɱ���R�S����?W8�I( �ߗ��'���N���ar��A�O�#A& ��S^|(�JG�:�A�Z�g���ȫa/E���o��7��F��
:$�fɾP����Rݯ�� ?��-RU�#v.?�E�𓑘�>�U��������!2�B���?�?g�:֟p�j�����:�c]I׽Z�;ɘ���ƩW`j
��\1C:b�:�y��gFAi^�h�X�_����FJq�(�*�^��%B��/z���r-���ޅ�}|�BfUw��i��x�Š�
�����y�9�)��h���.�7�}��>�瞶��e)�f8>�H{�����R&@�
e�lC^䗥f���2"�sg�2P�1�M�82�󉺆mALc%{-�s�3�|��5�>z����w[��4	����n��0��Gn�s/�a�?@�^&��O�����V�)u��F���)����P�:�)�!P�'^�s]b�[�m0)tZOW@>N�r}(	KE/�7OX䭾�s,�NaJ*�,|g���7&Z?b}��:��8��ŋ���8Z,��B�����]����z7�+i� ��O�Q>8ү��/�Q��니�Iȕ�PJ�r��f䖟<(5:�f>�޸�a������!".����}r��d'���F��;�R��֠q��-[��/��{��QrwҨ𻊫̬_�j����A�^:a�aYy������$ܧ���:��M�5�Ӂ6���R��bV���[{���Z��wFb�2��GN}ܸ~l����OnQ�T���(@�h4��j���[���z��mCo'i�V��[z����ߣ�����[s��n˄�LE2�k�1p!$��=����T��]5'���O��w뻖��X� E�ز�����D:��l�j0�f� ��~�[]V2��<�����%X����x��dO&+4����ǠR�O��3�qͰZ1jC+���/�{!m,k���ZƦP���~�.N�6t&\Obd�qh�0�Yr��꨾�[�Zᘘ5���O*Oa��������+x�}Ӳ���oYՈK���"�YF;�$-���
w�V]�y�K�\���<,� 4��b8�����rDa�f
�#�� j��!q?xe ��.Gy0��p?.
���!S\��@1�v̇P�9������QC�U����A��!{B�+ |������T���\��Q9�(+�@Q�r�N⅒��vH}��Ξ]"7�IZB-�Q�k��tM�$w)�l$�
A=|�D�!�a��O ��M�nq�s��V�-{����i����߄}䥒DP�L���_��@ߋ�V�,�?���T�ZNm��� _0�f9D⊵��~�O���b��kD$�z�k:5d~#��Rf��<��	�쫌7�&��*b�.��;�c�+%J���lů����k�M\�*l)���2P��׭%��+�*��9�����"�;�&��9h�A����'e�L�'����&�$�w��)|}ңJO0 �ʩ�2�W��&��!fUjƩ��v��-6eҏ�.>�b�G���O����%l���e���7�>o��HۓGM�r����!C�E��1���b�_��Zo#��(8��*��Re�W�Oa����e�w��{��	*�T�wy�����YO�,b��K�o�p?SS\���@Ӈe�M�`��Y�g��ݥ��W�k�G�^��[I�+��Q��$�ȭf�Q<7[�Q�`~<��	�&A���Abi�p�},7�R�%�,����O��p墯�΄Fd0��CFP�f��3(�5��P[���}�q=�vl���hS�rP�~��w۾=��'�:�� P�,��m�L$��;��y �u��]A�\�B9F����sMIF�
/I��*�����\R���_������@ʯoX��0�ة7�q���ͥ>9h��O�<Iؓ)~(�Jޅ2y9/Y�_NI$̃����X�0U�w�HNC&���f"�z��5/��5^�� ��G���~>�_��hdԈ�çF��Ґ���Wh,�ƍo�]Ƨp[�v&��]��'��Y�O��L_p�(H��9��逩[{ ��� ňA�jG\X-	�+�QE�侐�8�!� �������m�GX�Pf��U��{]�^CP�?�����R��i��U=�U����~9µb �`�� ��"��(<g�_}U���l�Y~������&O1!(�S
7�Ǌ��R{ɛv��pT�;�s�����0�\�v�'�/8�@CuTy�Bg�����oo�]y���ƪ\gB�&�U�`����xa�o<�ۉ��T�ŧ�q����ì�C����5���Z}(I��5P��yldݟ��"o�Ͻ���@�'��(�@`�pe�{���ϧ���� �Rh��JQnbO^p�Hi�ɓ��2�oo ��|&�Jż���$�R��n5��AwM���u(�جR$"�
 Ac[sT����7�,��pʇ��tb�+Ɨ�٥)����C	��R֤&$�6g��#���p	����r���H۶�W�� �6����i��-].57	�m�MlP���U<H
�[�A�gf��B���ER��4.y��t�ɘ47'�l��1/���O* �1G�ݾ�����~���$?�[�M��D~u�R�
8h~�?4G�K%R7�E���}�N��p7�g����;�����mFy/sN$d໌�a�׉�Q�q�_�r���벭n�Ķ���j,�;���$%�m���h�ǟ1�=g<޻����L�+a.�V˧a�^�]�w�"8>�8\�ZU�X:���Is��^�e׋P��W�E�}�|�3�{1�$m;�q����\�:i�2$P]�[�\��k�X�Ѷ��56�N�C�0��;��0܈i��o���}x&2j_�skt�NoP,�����P�*ƋH��f����}�m(�:o�t6H�I�p�b!�E�����c{оu!�,t^k��W_���bjY8�d�b�����+_s �*̟gAi���+�Φ��/�V�����`s�>ݹ.{�Hs��q5�;G�͹�-]:3g����cwD[�y�ԴܥRb�U��H ���jo���V0� ���ƌ �$A�I��Z)	QO�S��=fCP�Ҧ�=��KPf�����O
����̅�&��i`�B�<tLX^��؎��6$�B@ힽ��.���/fpY��,R<(1 �1��R���q������ s5�����J$b��nl��~��N�V����$aL���%��52�K.4�+_#�onMOK\�R�D峒kdUB�U|A�w	�9�>�.�zł%Q��>�n	��N�4@ܝ�9?ypsZ]0���Dʗ��K���L)�d3�WT�� �	A?I��9��r��n�x�E$�h��pf��p��vO6��t-��o(x]D��b�*H����:���4�И*������<�Ѷ|�9И�;8'v�xHω͞��޺jR!���-�Ѝ�8b��'���'߼�E!��ڔ��/����^�ǵ>$M�³-�t��ZZ��@.�L�O!�x���P��Kʊ�BR��l��H
��U*��c�,��V0>U=Hy�-�94!�� �<�|��P!U̴=5.�'��ȭ��=�=oR֯��A;�a>,��Y�h7��q�V�ד�Oar�֜��;seD�2�[]5�/����ݼ�0�H�aX!8�� �E}�'.Y�;���/���:��(N������!ֹVkD��=�m*~�_�XH���in�PCd�޽��˳�n�
�	��f�h���b�� 3#�Q`�kD�)��a��pE�����6^�c̲�K��-������Cex�V*}}Z�c��Q�f=�W~oE��9���tBcbg7Y���08�겣�ԅ1������E�L����˯�H>��/yb��X5�[������q#��H��P�T�U�����\Z|����B-7-`���L�&�Z�������-�m}X�̾Q�oFU�5�j��	�:�	�)��{}G�!����	�jZ`�x>�]�Iۼ\3-�|�+�p�+��8��� a�H����R���Ģ�]X��-QAraE�P������0p7��.����M�r�-����P��=��)ɠf����� ��#5���;��9����w�����\�2q��<��4�)fi�����E�?����s��
�}����q}fy���wiR�H�j�]C��\V��d���H	ȁ�-�U�8lm�Whxǰ9}-a0���#zFJbVr����E
��Zs2������*۟UCà1|Q�?�6��7�2�/mu)U����42�;�}�I�w*�q3!�'��Wr�MWOUh���"͍ծ\?���E�#U��3�'7?D����@$���(�~逇S_y��x��D�y��^�����r�Zt�|F	�='U�}~�\a��6Y����Z��.��:t'�BԄ2�Iׄ3���H������+g�P�v,�F−�;�:��n�h�6f��vb�n#�� �=r<Z�
z n�R��["�ǎ1n�Yۃl4��u�i����m}�K6 �ɡ�re� �ͻ�_�o�!��i���`�F��,�5	������/b����+*�~��e|�5j�O��c)e��Evbd�/N`vc}��q��pK�3SW��^q��A#ކhO�zH�8�NWks����`����f��n�)�ˊ�?�N�p�3�j�9�:X3v�uw9L:�� �c���f�)�he�}��T�ķ�^�n�!��'��v?sSN�8K;L����t�2F�~��ϸ/�4�챘n,9��~d�?^�4h�?��O����������a���HNW�.4u���"���,t�����{�?�	fW���m���� �5���yC�/�B� �`�N�����*��<�1?�G":Db(�?*�Ӛ�Z�3b�Nt����W���}���ī���$�����>���֜�L��F��@1� Zd�`�%�ŘT��}H��t��Y�\�F��_�̿k�j�����J}�R%r߇���| ԖT4;�g�#��u��Z81C¢b|8���X|�� ^��ї��ER���`�9��%!�Ж�`L����+��@l�~�-�����������[��'���G�����pm�t��c��q8eԚ����$=�� �����W���KC�4�Cq4���G�<+w/�f��X���+���̯�F�i�!�շ[�2 �����>Wt�|�"LZ��o]cȢd��9$�)i�MI\5[���sb̹�!%m�S����?/!GW���C�q.�� �g¥���Kxک��8�r8-Q4��o�����	>Z�?o_�&�lm _����\��K�dv���c�j�:�|Py|5E��2c��u� ۨ">v!��x"���a�teW�`3=�-�����/�D.~k���1Z�"'�nF3�-���^��ڡ����u��Auk��m�0�3x�w�q��Z�\񘡇��D ����n��I�갢�;�i�y'�$��p���y��f �I74�F�o�G�!��� ��gx�\1ӣ�G<N�P������H��\�;Oz�Sq}<�,+�\�W��7gF^��ֳ�.��9-����re��rj�k�� ���ه��E��H|�K��uUa����`��K(f(�P����N��9ֹ�).�Z�Qŕ���E�[���m��s�u��֙~0C=5��v>���L��&sB��O/��&$�*R���8��y��A���@N��?��>�&�oɷ�!1c��7xFE�� �Z������8=�C�ZOa�?�_��Я�;A,�
(�T,u#U\���V.�:������x�ac�N >Yx��!��q�y���"v7Y��C���̐(#\n�0��*I�o�s/3�*�y0�h�S��4�[���C�Ӣ�(���/����Hx��oؿ�/P·�������A��F*�.#������9�O�~C! .����A
F��}���D��ԟ���0F&����Z�՘E�>f�T�д�z�i�5��Qx`�þ,�)Y���t�bB�'��b��_�aCX�"�0�:�H�^����z�L&��N~�[Ƚ���Q³o)�9ڱS�?��[m��ZPa�P�Y�2���V��{��������:�L�	��4@bU⛤��S�O���adeFF}wr��\�3ii�u6�@���t)�=ѱh_&���k�)��S���9���v���S����i���PrݓU��v�i�$�_r��V�L��ͫ�##:&%�Eh:���x	��1�;~]�'I�p6@J �O.h. ���.�H�:���D���T�����%��>�q~�2��Mf�6���S<���3�9�=�؉��~�U!�x�M���Op�I�Z:C�M;��HQ����x���V)�����F�s���O���#�����`R2���qyT�ݯ��]�'�����)�`ey�C��t� �� K�7�2=k��fڀ1�'B���n�X]ц�E�Q���*�,V�*01���}��[F��u��E<��Ǯ"��,��zDx
H�n��w�\�J�w`۴I?A��3�8c�"��J��+դ��w$<�_0��=��!��@^�Y�������������Y��
m"�?���#���ͦ[B��ڢ@Y��������L�	j����+4�ZM����[娚�܇q��k~������ɢ����$T'�&��0ԑ57��~���S�YM����e�̖RD���`��B�0�|4�����H��9}���0TY�y�������o��X&X_6�Yp.�[����TU�ʷrl
�Bd����C�<���ӟgb��Z�1��b�-C7M��H!y���E�b�����*M�?���)�q�K^+7W!h��a��z�ni�{�����¸=��:qLy�{�9'� �[�k*�I���2�cyi����w-٣?t�0�-�^!%�]̻b�(�{G�y��|��G��M��x��*_�Q�3�8�;M������[�\�o��D�G�v�����I�3&��0�9����7�#����i��5��ǂ�R�8W���V�ᖒ[�p�p�^cq��������L���B��s�=�HX[7%�Z\�>>���0��6)|��|j��f��E�E��N �H��X]4��"���釉��Zx_^r�Q���Bk�C�����o}f����u*P��j.e�_�$f���|B�A�����[��p�D��9mQn���pw�8�3�D�B�����8�3۶����Z���思4�0P�(�
)��_�q��5@��;�|�~-]����~}���)���# Z�m����&������f����,��'��t��7��a�ׄq-;�"���Jr�A[��PJ�h�<I��^��ur�6?��H�M�	z~�D�ubZxL�ݴP6���ҽ��=�D&�v7�s�}�H�0�X1�F��C6	�5�{	㶾�F�ǖX�k��(B:��D�'$��LƜf��V��n�6�e�����J��{N?�c5j�qZ�<�0�k�lޅ���U*m�����y��HKA�D�:%WGù��^5�S#�ѓ���]���k9)�h����_��,(�Z��W���"
���R;�l��?��8��C��k_�Nl�}�pc�F�]l�§�_>�����Sx���3��R��E��|���z7K��J���h�HoZ#���Ŧ���J��Yܚ�HBj���fyh��'��ۛ�D��NM�?yX���������/�>�����|y۬`)���MF��B���5o�W����I�ُ���h��8��&C7�h���'z�,FbϮ/��A�,`q�1k7�^�3;	��ϑ	n���좸�[jur��C��?(����l� 1��ʌs|�ǆ��4���t�t���E�>��[w��>~!���m��cPpȠ&�iG������VB9��"�@�vPjf�M���C!���u�민 �m,�嬌���Gq�j��F5�����@9>q,�m�zT�iy
 �<�E����w�/��X����lY����d�(�9���W8���&n�&��G˧p4}��n�l���w$0�2?�^q��@��.�]X��|�I�3� ������A�.����J-Љ�,����M�8<w�q����Mb{L�4xP�8�"eO��`��Y���߷�1+.7�
�Ը���ݎ\ud��h�9��饲c`���YhLW�uu�\5o��.�N�����m��y�T���S����.�/�qn�4�Yo��q�&���H�+	y�2�a� L&�yh��eZ��*�����w�
��7ZH ��&C5�ff�7yX�}�X�A��#�f�����a\�����PƮ���`A�h��@�	�R��1� lK5�vK4�$\}�����r��Fs_ɫ��E?+L�u%�F��+��j�~ğ{�M9��W�{������1��?�d�BEb�g����U�s�+�#d` Zw���t�X��W��"��J�8���-�^=��XI��:���oo~��*����Q9�(dN-U���t�G��y{���1^~�E5�5�f[#m�.��?�ؼ�+����"�:���
�l�8��X�h-�%��S��t0kh���]���_h�Ro�\3���|r���\�IDΏ�ᖢx��x��Ll��:А@�b�$������=�+�lR��w�������Z��6���A[�^�ٟ���#A�6��Sp�g��k�]��i9�I��Y(��Pل�U�9÷�,C�h+�6"��P�*#��A����+�ԴV����0�s���9��{Y��'p�X<� �U��I���2
��6�>��DTy�����y����Ԩ�)j�&���y	K�9р��&6�j�$9��o���M�-��/���y�v)��׬*�/ <���G�.t���8|E?�¢,�z�ɣgј�Y�4-�D���Isj%��~���w"6�4�Z0,��`!�%y塈Y�3��<[V�<�Cͻr�ϩ�dJ@J���3(��zѳǢ�R�{�՚��+��o�&�Q�:�W�ł|92�}��6�C��	S�)�.Q�����L;,&�w�76k �����g�|�tRy�&m�_�q�����ruQ�62R=��AXG<��~��r"�fϓO: C�B���J<
\�t�H0��3ک�;�x����@(���nI����cf�C�3C�M~1@_7�d�:r��T�����i�Hk���8�f[�_�_��X�y=��*���ܧ�(�~�	@� ynw�0O��`�μ4����a}T
aq�K��?��߇�΄|(�F���j�@Ӏ���*�T���Tk�m��5��=�t*Sdf��*��MC�������r�O���4���V�M� D�A8�~-�4�1&�1��}���|�O�����?o>�_�x��}Y��p����y�؃�P�g<�K�T�ȳ�K�M�g��n���L"B��=)u�7C�k�-z�=$��O�R,�Cf���u�R����D���60����s{�fgPj_7Ӽ@�#'����]�َ�Ь���G�	�I�qu��9�G���t�l�0d��*
]8�,��L� 9���ⵕ���U����A�Mm��֭�Vbfz��@po��� %��AG�,pE�!~��P��lp�h/G�*��)�����/���A7��u�J�ǅi�;��)[C����'�Ďd{%�SP8s������9@��w�w-��}�����c��54?���[V��IK�N��)�4�·���}��y���f
������u5`O8c�m�at�0�@�v�=«M���ie��Tr��O���|p�����[��Ŋ�ݫ���Ed�G늇����%xTQP)���\�����r�(W`���~��ʫ���䪓(�����P^��O����\�$ʧ7���>e��$�-L�h�V�k�!4�i<+15�}E�[��Q�ɓ��u��__jl]��^xPh���smv���k$�[L�;!V�iv�w�d#�)!#_+�adHu��l��k:�*���r�:~�&������=$�s�j��sIe������H�h��oQ2�f	
<���"��oߥ�҅�{fU):k"�&�RGD���o�'D�~O��Z%u�U؊���l��`n��!�0'u�ګ�i+ & �\��ḱ�/@0|2�j�W�s�������T��_3vQ �v5�B˔b�x�Q-
Vt����,�*8��!��}�`�1��.��x��%_J,�%&���� kXqR<)��°�A�T�!�,�ى����\p����� VG�Ƹ�O��1\�������2�g��:�_	Sv('p�*c�[,B��.P�gT3�/7��W�v,�S=�f���#A[#��;��Oъ�����j.z��A�=1�d2��x�ٱg�b���c�=��~��R{*�{�ߵ���漳ʢm�{���������e�֡��C ����R���\��d�`a�*)z%d�bZ�^�-!`�T�jo�+���y�Kd�>�ml�p�!�SmY�?	c7�$�+{��BaWEФtI�՟���Se�s������w�B��Mq���Ȝx4#��=.r� ��y��s��#��e�(�v(]�f�&��7.��1�O���l�"~͎��
�d�I'��W��/Wy��w�Ap���?�_o��2F�nN�j�7��H�t�5�X|S�/ A�lb=A�+0�
�] _��h���k�<��w�~�#+�N��ܬ`��D�|,���V�-5�=6U�,���r��造����0v�T�;���"��վ?����uq�s,tmJJ��E�� ��S�)O2�m�l�j�Gw������Y��>�;�P��~}�T�5di��>R��b�w���M3�Ƥ�I�p�&����-X&焭+����2B�jwC��:?��kw�,�O������#���Uô!�ۃ��3�Y�W7�K �>I�]�ߌ��)�u�q��	)_5n2r�Ֆ��o\k4�W��[N���>�;��E�9�)��U���W�WoAJ���k��Q�5Ɯ�4s�����e�_�u��_��������N9t�p����,1�1�n��D�qn"�Ɩ����Մ�,Y�>�VXT�%r�ڐ�)
\p�G�ο���I��@�����˨����0��߇'D�@���]�mѫ�}�,���U���!=����	�bl1/�+�#�O,�[����@��i�n0�>�W�b��.�nS���p�K�P�;Ug:0._�6��]���e��V�Pv�(���~��^|���7�2�X%���K�z�ye{��Ġ��H���$��_�p����s���x0�̓�|v��}�@�@%���\�L!�.��^��,<��(��kK����2��,=U�Tx� ~��$��&�Qd��R�����W7V=���Vݙ����%/7H��	 ���mQ���7��"늖ΰa�o��G�W�hߥ�.S�JP��G2:k��;09���R�F�= z���B��F��6�z�tz]�`z��t'�(�!q�����%(�5V#-�E֛��a��It	�U{Dp�;#}�`C�x����weV��\'t]H�7ވ�$����k��v�i�%��!zW���BW�;�*Jzn-A�+Ď,m����l@���B��e���
K>]r(
5;m��n_�������[k FSK��5$��XTj�0��ǋ;��]�c�R����	�u���/��.��剛�Yǌ�J}��j���(~��ܖ����Fﯩ��<�*�6��m*V
�')�	.���aD�N�0�W$^�CG�_�=�7rt���Lbr�1"`�4�̄J�n�ǽ�E5k���l9h!:�N��m��z��Q2F��Y���Y���Yo֚�)z^���{P�y�AZ4�쬈��p������FP�A-�>���������/��О���bT s����?B�?��Z#I���D�m� �%OzI�.�W�
/HT��=�9�0��{�ݮ�-���G�^+] &�� ЯF"p�����a�'{�N8{�����)8���\N���w=fzρ�!�h�0E�a*�|�M�Ho�(U�:�#�4�3d��9(B����o���"U�rO)� �fl
�Z�)M��J4��O�}ذv`�MV�巸��^G�� \� ��^�������JZF�v��!"[Gw���!����ʪ�*"&`����E����8��FK�y��}�z��6�8�ROc�Gv�* �r���#���@���x�A����K�h���9��c��>��;�� Х JF]TK��J���T�j�C �%�q��}��E��x�ş:k�-G��*~��E��ܞ�噰ɞq��}�q���%�M��jb���}g�!K<�a��7J�`��	�ѭ]�>�ڏ'�.�x�z�Gq5	�#��y�E&�(����'W!jX�0a�!_�H�bC�Mn�V^P�f���W��!t�,����pmd��;E�<,�{������<ؚ���,�"����oO{��ju3�۱�=�ٹې+�@T�w&e���lb�8r+tI����}2�\�����\�@Y�.�&4�'������p�/>jV��;�����Q�#�yD�'���*0b���5�<QhG_q� ����l��Z��Ϫ�鰛�e(�����$����0�� ���V���y˹����ҲoSg՘vH����^6{" �����7�L$�vE>6:5�?�_p�US�jKm��Q2~M���u���?�Pբ��^Yw�Q���[�-�]�W�����-�������uX*�w#n���5���w8���<�5����bC�l��P�a��&3����'M���5�n�;U{�X�A��Ꮌ��k�%��H��2��-22�丸�h���j�7^gG2myO��3��O�L.��2�֘!��`���ܵ�*�`�Lw�ԗ������J&3~h��PR�����n�rV�K�o�1�`�'u*�� =7��Oc�<q��kW�WM4����e{�P�a�pGn/5���P�3_�<1�)ߩ��Ɓ�u���_xm֒�_�	�P��T���4��ʏ���-��X�����@��%FB����+p%��}ajM"'2���0�?���m�s�H��?_�i�����p8�Hf�5� Eӽr���3Zt�M7�l%�q��CJIW�#�qcY&�M9o ��Eփ�`�	�:u�U�~��
�5����TGIPB0�:�����6,�cX:��aQ?�a��z��l��b]-
5��M��0�r������=�U��l!P`ܣ�9P�kҍ=�_��oN�p�2�2#��q��lс��@�b��&���]Ѕ���$c�E\��3�����0,��@��<�ė�W�;ӳ R �lq
&�N,$�1�J%�N���~;��h�h5��]�=э梋�KZ�� ��RbZ(�h�p�����$�g�#�6'�w�O�  �1�Mu��Q	�D�'8!�찂p����qe���'4b��;�4E�	Hղ�G��<����lR|�0A� DQ��*�l^��TY��Ò�o�w�ќ+O��Dl$�K�kJ��6��O�*.#�O���4���S�EC���P�J8� ����Q�9��t��o*�$��j���BW?���&��m	����R���ή�R	�Ƒ�h+���B�zK��qY�k�'�F0����>H63��Y�VY q�)�)�����I!d�uS6'5?��n8�bi@�ܺ���:x"A�Q9�s�sS���P��"H�<`�K����4ʏ�����e!��Q�}9��U�iF��¹�2��ۍ��ћ�*�m����v��
Jf�x�$?c���F�<Eh�y<����;L��3Ó����ǞeF�"(�Ho_�;��|�_��~"f�D~�H�� ]	�p�s��w1B S�.	�7��<'����mت��(���CX�lj��1�i�XL��	;�
��BrS�PZ�b�aR:~�J�*#,/��I��o��y.�b�kfe�0|�Aph%]u (��`�q������9��:~��Y#�����B�x2w俾;;h���t6����|��T-�
���*��f���j�{TgB;J��7J�&K��a����Xn�5^C�Z�!=��h�U��q�Ȇ�Ѻkj�ǍЖ�Ґ��	[��\۱�3x
��t3�+��F���e�"��|�E/���#j`5huG�_�Z����b�ں�{iMEw��Um1�M<6��]��x�@���U�ӛ���#fT�����ɆlM*4�Ռ�n�\�-Ҹ��@"��zJշ~�`�H�G	�3 ��:�_� ����S@�hl�qV*�-Gw�:+`�ˀ��=��~ȰRGr)�2>���m�?Yhff�{�mj	SkB�\�+$YjЅ�+��/S��>?�8��@�l�����$���T0w���"�H�謪���@��<u����m�<>N�.&���g]�%X��`�τ�Ǡfq��骭i����
CQ؈�.����`��61��D�t�'�����v�Q'�5�w*w�sV_���Y�M�t���#���fa���n�� �������V���R���%�����ʘR�S!d��*#ЎgzV$Ltٱ=����w-
ܛ\e� �e����vi��򀵙쿆�^~��`�e;��J`��ʐP^w�#�y):3#�2�8|<��-��ŭ�`w�Ĵ�F&���͉DK��Py��j-��{����Ϟ�d|z9�������r�	�
�dlS��R��DI�����V~n�?}Ԅ9��"�Md[��C��D}�d7��}����V��n��_�>�)�3���E0�r��Y�T7i�L~t�������n�۞en/$Q�T���Xk65л�b#��@8$��}Veo���g}j�Ǔ`i��}���nf���`EH�kBܰ8k�޺gy�Ϣi5�!`��0�)�Į%��)�����@h,���U����kc�r�^~5�I=t��K�qi٭Vp�g��!hI�QY �b���{�#� K��o��H�Ln��EX�]�+��F��ԳИ�3���B;)��rK�(�LVɽ]���A^lX>1}к6���}.4VG�)9���Z�tRc�ԃ��s�uȟ��)�`��6�K�f�����Pᢎ���?�3]��J�}g���s�&�$>�:I���N"�(�(%� -�;��Txu��K�o�D	���6Ų��>��w�_�Bc8���-`�8�\�U(a�WB~�6Fc��X�	~`�G��'�-FS?/�L�R׹
��c�`��#��W��rRT�$֣�d_�͛��t��a��j��b=�����`K�8�}�qf]g"�|�/=�Y��z��H�i�z��l��ٿʤ��-E������|�T��F,���L偖l-4"s/�cW�OAu-�r�%��a��"J\�wx�h�Qj6w�*vG׫.B����gj*�C:�����*2G�������l�H6����S)��U��=�$AØQH?�Xދ�3�������0A3_"l9�*��[*%�[��XH� �=K�.�;�9�J�d�aȞ�59�wA�.��p�f����R<��d�佊]wq���OZk���`G%�E*l�^i�M�f�"D����
�N�r�TW[���v���
��}>�H�|�WDM�@����*3�]̾4���y�_s����q�t�Mگ�Gaϵ�9���6l��K��a25u"9r���t1HW��Nю�Ey��uᖢYnVnuM>��:%����Ck����ϸ�<��=(��<��l4��Bɳ�_)Uf"�4"p�[�B�Q�=��%`��+�����52�U�B F.-�!2Ye@��c�
�d�e*j&��U�q>�~c=3%AU�/��EwĪq�_q�C5�j,8|ϵ�N~^`$|�m�Ϛ:#�.7�A"PFp�$;!p����4���>կ�����k������jI^�!������:���u�lz�(|�ͻ��g��;���?���L��l�ns�)RTD_���ł��X{9JEF Hu��z�S�G=2L2en�	��|�9�Z<w��3��S�����H�l�����k����(2��dI�B��Z�R*�b�>Q��D�=e�4W��
I�9h.f���	�UJ*��CCL��5��S�8�ڍ�Pџ,�~#���u�����ң��Q!���)�J�.��̹�yK�)���a3'qD}S+eϊ���&�� ���b��e�����R��}y��3Xn��%�QX4V�C�{��-޽#X�����H���*#gf��9h��y/C�s N&�;��FMu;=��F�^4G�C#G�@��	�L��������Iq��fjO~��׹eK_H��;�~�A'���ĐJ�^^�tpj I^H�|���C�5"�mG�&)��� #a��Ro�g9�G�_FJ��H4��0�o��J�;w?is�@���D˿O���L5���lI�m����>�*��$�V��+���XӸ\���Z ;(mP�ꥦl5�cpyY��h�o[N��c�T�{PS�Q�5|e�q2�L�7�k�� U��ka���}��� � e<ɀ喿U����5a�~"���J:�o�c��­���yaI�����ǃw�zɾ)��-~xüd��R���j�"���|�Rȟ_c����[|�w�����Q!�@�i�^G�hh���L;�*��WG��/>*`��x���#�gR��	��Ԛ�V����ӷ�fK��EE��qՈ�X�g���<ƥ��E�E������3a6;��[-5� !�?��N�B��g	1Պe$/F�c]�Wi���U�)s�V72X't�̊3��>�u�XL{z<��)����HC������A�u�l :��Xuq~?��A^����h�����7��ٙJtb�1"�]��x���ۜ�z������L�O�����\G�.�Xޕ�AhJt�D�[�W�m����	<g�)C���D��'�2/{��H��n)8�J������1P�5\�o���o@	������_ڵ�H�a�&��R�@c�'G�
p�fQs���6
��5A��`#%��{����hsU��X��G��FQϹ>H�t[~�7�O�u�[�  ^#���[,��(�U�,��+�0󙧆��n<f\��n�*����rexf�&��b`.s�؁��j5�	%G�M���p��=X�����3�
I`��jkr���)`WE��t<g����Y�?�j��9�$�E���LG����D,zO�h �qI���SW2�z��z��*ic�42��k�	C�����kʬJ�/c�΃1t����=���B1�G'r�";����d�iI�n���n�;kD���@����+G��S�=�V0�TD&��.@�VT��H��(����M�9=��T���?v
�(����'�0�\�[���y�q(�R\��^�!EA緦�.xh�ק/m�q���RR3�T\�a����9�D��#��Eϳ\��3PJ�t�Xɾ?m�z]���-��ڝ��}ٙ��U�2m�P��Y���f��Ʉ�����Ɖ�~Nd40:4��6��|�������Sד�o`Z˄W2�i���!Һ�o	�_�m}�϶��33�Hoa~�LzUҋ�z��[\�r�����a�C�W��!��,qW��&����	 8��[�i���%�r�~��
���^#p����`���Lͻي�$�V&*�Lp��\.9)��-���>�X�:�HD����/���a��z�˴Ɂ������!��}�0S�� aܠ�
�h����Ǿ��pNKm����XV)�_]Ϗy���Q7ι�)��MDc6��#�~z{~�����4��c1K'j���.ڶ�QS��'/�n�$���Q\�]��L2�Pq�x���/�σ����J����BOgW_@B}W|�5�9e�%��7o-yy�1��q���S=�>�D�m�Ƨ=��RU���B���=س�0`ʊ�cOŒ<R�~�ݱ�_贕�bs�e�]�FS�j�����&�Sl��ߞ��i>��$ �g���	���#i_:��x���c@�4)!���]pRl��g�����2��͠$uF��P��	������� �X/.��M9(5������R���e2��H?�� j���<�n���1��cƌ��:e7]i���2rx"	���Kj���(�BJyk���R"��*f,���{R����c]0ߗ勌�pf��a�κP���| ���N�P��B|wR��oH�R:�E�E��7��v<���-nJ��d��l��/��t�@���O��W�H���~�f�5H� #�Z�>��'I{y.tl��WЎ�'��co��.�� �i^L;���+�ޭ��K̟~�%0�d>�j�Z`�0�X������m1�pn�:)�_�9Q8,4���讁����6�{��y����J:V���l�VB�����[���7�J.����:�^��t|��ؼ@.z��"�Qu4�ң����b��}_Lz�RDLhC��q%�)q���fGzz������+T�D�D.*]|J�l#���9�[�̢�����zSx缊&k���ot�擽���{�����!��J�	Ҟ#ρ�b�N�]6 ̰Z<fYw�wH�B��(�xԜQ��j*��g��w}/��n7t�3���0�/�M��=�ZBǧ��8�Dx!*E\q���T�9�L�h�q��w=��9��?��8{�^q�e껏e�5��<�ڈ�����`�[�-B^�(�9�\L!��'��}�ָ��O��oc,���<�Gn��)TZim0�sQ��O��+�"Hֱ�v�^N^�;���D���?(M똲�Y2n�&r`�������#n�7�}�C��`�TA���ڶ�q:QW-����M�:_��2~�eJ8�U@��IX<��s��
��ra��խ���P����vC����������ѕx�!�unI�z��{pV�U�a�|L\X��g�Mm5x���K�9R�ќ�f�6�Gh��&�{�V�����
b��/f���*"�D��H���K�!��5���	�djN�Y<L�������k84"�4����e  ����%��(���Vhgf�l'l�u��UnxP�������L�
=����?I5b��?^�#gD��g�Q�@3�]�Sn���/x�7�#�3~~��s4;vw�|��kݼ�PnHI3�A ��@����*���YcL ��U0�ʷ6�������,����v��l,��دh��-�M���(�\�:.a��W��{��6�]����;5����	�m�ؔ� �[7!�e;�����Ë"z�&iW{�&!;*�*��Z�Sfn֚G�+�h)��6��8�݅fu%����4۟��'놮/eOp�x�*�^�W����:u��d!�8�$9��\�_��UP�����'݊<6�j�h,����'n��Z��w-���QH�&��bgcs������/��R����˾���giC7S)�@����w�Y��`bģ�<�U�%/�	��T����%XY�Ei�ǩ�҅snN�Y�J�2��|�����0#�	�}]���I�A��	q���ο:%z�m3kJ����Ɉ�Et���D��v4_��B�w��?�Vb�w�YK��%"�,L�qM�f�W���P��|xt���z2�S���Q���-�`�x�\���Q��A�2�@�<���M��X56�[�z��*ղKF?Q�_��pO�ءu'��L,^�['�M�
��ɫt��?�`B�4�����V�S8�� -x�)��;�����v9��D��v��>P��>2h�nkz����3Qzķ�qQC�uSM:��ak0�zwaą�F���%��m�P
����&2�l|��RjW���Q�{}�drw�u޲X���^�����-~q�q�� 0��e��Ʃ%p�/�-t��B'u1)'�,�_�ӊ��C�54#e�ؕ�߻�*qiыG�p��5���A��fj&�j.8`�"M"V�62��ҝ2?T��6���=Fq$Ւ�k�z�B��(!~�̝�w�$��m���l�؅�������#H���Tn��v<
��
 ��Y��/��Pl�1�Μ����KiS�#K��E�6�{�@L_]�n3@�>�瘆����ԙ��!hX��AB(l��)rEh{���2[ˌP(I&
�e�.���~2���x��c~^1*ᯂ��q��q�����j@���7���Z>�@5A�r��kȇ�]�nWP-��cKq�X#+�J��H�q�\���!��Y����jf���ӪW��#hj�W7P��H&�@���gQ=_�e�9:��Ih��Q����_��<���� �4�Kdj�xOD֧��E!��	'ׂ�ɑX��p(^��}p6h�7R ��������>�6���M��ɿTlb���C����k}Y��@�9I���q�<q���2�%� �ċ�i�Ike�"��7�E�l���k
\Iu�>��4�#����:w=+���h���4��[mNjC� ����'q��'n9m�Rd�5R�W�.;�K��;�`O����)X�>�'f1H#�Kҳ�� Ɣ
����o�}w��|�p6���)�I'�<]-;ͩ�du!J�U=bQ��l��F�y40��$�
�~������ط�J�����[��z��]�����������U���-�E���hE*IU�բ�	���f���#���^8*��6q "����B���ݿW�1�*����:�7���܉�$��@�K�dv��S���2��]Yν��ڪ����:��w5�1�eėa��kr�y١�67XƯ�.��"�{�P��A��Ă��#���*��HT}��S�ۆf���D�¯��-	_��X"�ƫ�\ҭ��c8q�M,p% ���C	Oh������n�[����R X�l��$O�jƇ��E�+F�*�������J�5��a�|�����-���Ұ�*���!��+�!N��0��檯�����1�!�{M�fG�^�-�0&�;I���k��������nj~������^�#pE�d���Ŵ���t�`���2��2�fǌ!RjUC�+������-�uba�6[A��YO�<�#���
p�z(������n�F��%y��$��t|�ԥB�i65�{���!PE���J}�)_kլ���3XP�%8��R���X;�6�Z�9k�w���	;_6o��S{@�u`p�V�\�=B�C���� ��T��a���C,�$�:�Ih{��te�\݀
ecn���y��	�rq���v�7���r�'1��������J��Y1	:��hWl*v���	���s�R=�bj�N
�W!�1Yꉧ��/�1�]U����N���1�2�瞝�[�[�y<��Օ���~���OO��"�@H|�ԔO�a{ I��I?�W�BVֱ�=l&�N�����+���+���Ɩ�;K:N�j�1({��B��~������g��5��A�!�_��B,��7���M�jZ�=���f�1��[��_V���x������/������,&4Z�;~�1�Pmk�.��S� �)��[f!�Q�_U'@�s�Ȼ[�_=�%U��ʺ�Ĉ����T�dׁ��j�ӱZJu�Mh�1���V����o�;��o���|Q�SnK-7�p�r�m�|P,�~��HZ�yۘl���<�$��w��$��ˉl��J�`�=p}?%�P�$�6��AĝB�*��Zv�-���v�R�`�k)ɖ��n�q)g��؟FCL�7�w ��Pq:�4m:��?	p�f���X5�g�Vcò݇����+h^~�,���c������ ��3�o���g10cOYƲ���h%`:9{�:�Q��#s���̷�ÚW��ҫ�G�4���s�=g*-fT��!��.!�Yܗ:TK�K��nN׺	7p� Ꟑ��G�6�����nnʵ6`!��[��T��y���|��q���Ҝ���R����T)�]3;����c�/�"udܯp\�[s�]Y�����i425e�5�\P��:a��9�隯O)A7'�h�R�$<L�w�*�*������X�s�P��~��������@�D%������������'�9�Y��XZ.�o� I��q�l���ף絗�Q��C���M�N�����4�ˋ.�
��p������@�lZv-���S';~y�>���ؕ�:��#�PK����o�JI"��v��]2�4ǌN��P�����a�{@�	�X���b�@5�TP�����r�����`�n���ά�*xZ�zS�SrOx%f�oݥBxe��s|s��p5�R�����,�H�̄�ИI��V�z!�洍��2����t^�y}�Ë��E`��w9z��O���hmWk��/�M/���y̟m�ʡ:�i�@m��k�	�T�+i�����F�JK@F�m����������,]��~�U� �%���N���*B�$%�����u0~��ұ��T�4B�X�ɏ����7��[�\>��T%�	~�끷�3������� ��<�{���ٳ��Q��^ ٍf�����lv�!(og�)�q��{=C[�G\�['8@u�͂sm�2��B��<��Q*�x!�����k4�e��d?���qob��%LmcT��p4?y���`�xSn)`9e��}�W����Dg|����Y��fT�;�'�v'8� ����� e�Q��m��Du��f,���}���(G2;���?���#��_�0&!$�Vz�*x�"�������/f c�+��d������5�T1�B^`�s�1%5b��ʖ��pk��f)��L�F���dY#�).c� *��ΫK���§�#��˱1���շ�/d�#�y��lln-�T���U��#!�����Ġ��%��D��J������;�I�Y2j@֬u-3���
��u�A"�ȿq�w# �b$�mޙ�����?���'.��C�N�'5�U�Q��`�kt̃y�!z��� 9_n���4a)�h	�&�O��o;���X�g�ٔ=�ݸ��+���+��(�([u��R���h����8L?J*��3�b�3H�!�1���pq�]%&%��B�N����P����3�|B��s�^ #��r��7�$v�مܡ�c�ތ���aX���1��{�ӗ��/�ku"ϳ�|�k`ق�_�y�7Y1 鸵Kҷ\� n��Ǆ�G[ԣ��{�L�A��-(�&B���:���Ȧ]۷V�>R���G5l�w�U~lZP:&|�zTU��*���zU�"���E!� �C��a��k�����m6�cY���e��]�f��-	޹&���=�ʩ��NkC�֯/r�y��㍝����M)Ox�0<YC���X�;`�6����#LLJ6���"��[X�C�U��|��/��W�k<ّ��bITp�ƴ���IsX�'KB��Bs�;�I�3�o"��ҘP���S~|N�b�AHV��e İQ=�cQ�$,�V���U������|:D �̕D�-���>�������@&�!�	8M����_Ȅ�-�f9@�c�{�*�pMH��3/0!;׵MlHOVA��U'C�\�M���|l^��;��{6���jR<��n ~fnLf��8*�a��!/�'���rh;b��K�'o�"��P�"�2]:6c0�<˼�����B�� ��|ߴ�92�M�c|=o$
����]��!���('�NY�l͎
ݡW~ȸ� r^�J��	�0�.��zN�a5��a�8�l�E�Z0
���H(����k15q_f�]m�SiV!~�k(b�y��\��$�7�>�\�����l[��p�'�2Ъ74���C�$��Ȯ�J���С�|i�x�!zx�����B��=��w_&(E#��j��uїÀ��Ù��(%pf�o����:��9������e�P�3��;�3��<{?i�Q\LHu���ʏ�x��:=	�zj���;<.��� *���^�<<,K�L^�^q��b_@e�YPd.�+M.<i�_���f��F+�Dz�X v��D�m� d���xMaq�('�����@86������:)��s+i`F�A:���}�������� T6���D�%��4G'���ߴ�F�Q�������'䕃#8 z���c>q�4B��'�P�ȝpօ����`vc��a��r:��l��@N �?M��o^P�ģ{��XP襉�=4◈�_Ž��8�'���^s9���A�R���=}�Ľ�k)X:��.�?N
u>�Zw
����&E�UL��Ĳ�^g�3��)���e�!��q����G�ɭ��8BǮ�UgA��_��p��l	�ڔ��H:0 �#ej9�"��T�`�mE&����G������.ڬ"L��Fc�q��\j��
5
5{�uXg9'�K�H�-�|�6k�H;zL�(�f_�y��#�z�Fů�OE�7�k����9�i5�Q�{<���%)�&5�ȖbNVU}9�����?���5�g�	�+�j쟼T��A��[�Xd�Y��YP�-�:�>�F�)���CK���z�4��������~򅱀�EM �58%��؋Qj�|��9uOSQ�!P��)6i]���/S�&�rH�J��-=��`���KE^�]���GWH�������6�Lz��#T���%�w5�x�[�`�T��m�󡆡��Nؚ4{4�^>�ж�1����'�W�Q9�F0�FeCO��y��g��G!�sA�PFG�Q(5���#q�e�S���Ae��}S� R����Cd,������0��Ӌ6��
.��!$�.��b`��;�o��a�)��U �����&�#����Ԣ�"��saS(�dN�9���=��̷xA�1���=�[�L��?��� S���w?|sy((Z�z#9G�N�ͺ�E�XKd��[��jm����4���v>����l2�b�.�����g�@�z_�d2-3���su�ų�p�g��e�XPᲸ�ď� �>+�s��*���ۼ�џ��ȟK$��L������g��_��`���V)rH�Mo�O%�HX�(��'�Iȝ���T��&�j���Tƕ�WN5q�o.�uEy	CK�VqQ�rr��&7��8��x���1�#d~����|G�@�m{ �8�w�?�����F�:X�
���!w�na����;1+�{�/�������̑R����[�nC7�	uȸ�]�w��#T4E����� k~Hpf�!m.��xpO��N��^�V5��g)�𧬲@Z�c��%4�zdЋW�SMi�2��1KIg�9S�c|CYME�7|�[F�.����r��
hͼP[�U �>s�ɏ Kc�Sh.5ګ������QhJ.��-\�u���Aw�A��&�_Y7�b�C��Q��
����\���[	o�(	��J�ʎ�2���B��b��$�p^?߭�rQ�u'���� �3p�n�ehMO��{R�4h���R����/�At3�k���%?��T6�jf��IS�²�Y�$Wwz+�F�6.
 ��O8G���m��H��������#H� ��đ�o�>�k�R�hO �`�jfS�	����#�;5S�M ����7�7�(2��H��P��*�_�=w�ƻ��q>�
�E�'4��k��J�w�w�Pym[Q�N}r��1�-|_���AR��b��n܈�D���{J`Х�aU(*m�Ŋ��7J�Xf��.��뗊�,S5����hs�O�2Ni[r�^��,�I�6ȆvG?�Ȁ���;�"���j��f�A\!n�ee�����6�+�G�<ma��M�څ�:ޙ�d���,�̗6��֏��nw�R�)V@�1�<��D@��\+�>�Y�
U@4?�t�_μ�#�Ht@�����Ӫ�9((����s�ԁZ!=�W�n}��˱��M�h^��%�
�%ʦ�ރ{׊�}.ȖmG��l_̀���!*��z>}&�}�%�u���.K�k<�=a2):.ߪ��.�uC���7`w�7�R�Q��F	N{�������+h�4���M��߯�C��Í�Ð�m�=P�1
�nÿ��|�#�G�Ut�榻@����h��`���_��K����x�����î�S��mb|P%�f+�_3�[���{�KVL�?�$)X5u�ɛ{gcI^%�!���I'��K#���ڰ~h��}��=��~v�&�#�I9��M�QF�Ͽ!�r��zU�	�B�5t�%W����^�	���S��f���%@��������}��
�$�D���ٽQ2jb�[� E�q�P������gAQ�P�o-�\����x��T��&Y?.����a�����0y]���~0�s�A�e=�H%l�[0�d>��$�FP��I�0��DHj9+�UZj��K��ѩ@�d�U�J%���#� p��$+�9�#K�:�X�pNʦNۘN_I��;��{��ƻC��!ա��DW"صp7YuxW�����r�e	�!!�mY 9�0dI�D���Ҩ.��i/D&u�ICMj3?:g�p�!3ӏ'��$��,�uu�y����Q�1�C�fT��3��F?G!��W�YWFC�Z�Ch�@NR^+b��[g��2��r+I�X�ȩ���[4c<'��R�N�|�s�j�g���o97��uN�fؖq�k�n�9�b�T[��i��@�[�ycӴU%>���r�Fu��L�p�s�31%�v���:��˜O���yZ�rM�˝>���0�H.|1��,��%�C	�}�\��N9����_ n��##jy��^E�V�Z�����-Ab�i�r�fmϳW��D'd���B��AI��2J���*Ե/ːg��'��O\K׆�BM��Ǧc�9�蝅">�W�&��]"z���O�� zp\T�u"2\�?-��y����]9�x���>u��_�l��#,%��E�z�#�g�i:�U8�j4��u��[���1tԂ���Ś��� �m�`�k����:�xP1֐�geWo�$�I���7q=n�	j�-�g��� oF�����5�LI�����,��ۦ4I翝�1�s����C�S�f�xȔ����~�;ۊ�b��;��"�:*Ǯ&Dr�����y��r�f��fUO�=�˽�����_7t���$�WKf�[9_���6����R+OPw���g`7�C7,h	�bD�����%�Q��5���uc��W�p;��K���n�	'Cg�V]:��F�{����t�Ŕ^ry㴧����h����;�|�EЋ}�*�oT�}��{�=o�������'r�0�&�am�B�m>f?V�]�	�R}zZ+*]Ѩ+�.@�?
9z w:j`�t����*L�t�W���CJ?۪���9�u��X�t�M3��:�LR�ֳ]��T�>����Ƅ�g��@=sˠ������4���{Bik�(��V3�v�<��"��|�0ȹSRa^�1��cr9
Q&�v x3���F���;��m�=�!G]-�2<툿y��J�ލM=ņ���il�:;L�@|_��,�Ö[�r��R��~�-�t_�@ɽ�;����hG_j�����rfPzV�zH��H6Nj�膾�|\~@q�D^�ʊ��(���7�� �?�g"k��`kK_j�0y�ēdlDBW�r��e�1���p)l"I�t�0Շ!\R�%����2��^��v6H|:ܥ���%�1#�J��k����V�����$��wS!����ǘ�c�?v�'+>=R^c:�B?��c�+,�;S��Ϊh��PZ�>;�ߝ
�hR�	���\%[�j��!�K�*5c`n���^O��4.�g]9�9:�?��P�d���LH����t��;�����k�K��'*ȹ2E�#Fj"�W��#�%|�^K����i�O��V;3���B(=X�_�.[3׃��`�*��s�L+wE8� ��p����x��jdd�RW���h�;��*]r�Q6@�*$X�H�>m�XK��	�	y�����^��FJ
��ci�TяʭA�����i�>7�� #؁��GMؘ�ߏ�]
D��|2���SBC<�k���`�ٵ�{#�{���N��h<륏���oSZ�#
ۿ�1&7�'uL�m����cU�R�8�}��تT�1?]G��i�3b��
_|���Ȍ�/���_}I��/����z�����F#n���6�L�
SR�UU�b�#�N���\�l�9m�p�c�Lұ^n��5T�X�
e�{�G���'sP��QR�ں�A�C<��V�_�1���Ǭf.�7�<Z�PwT5�;WJx��v�����Dr�B�Q��`��,�"f��qKi(8�^�6��T��_#��n��V��d̗p�)`��j�*�|8��p�!�zl��)b}����o؊�^x���|;��Ҭ�M�F�X�dѡT����ż^#(p:���J��8�e.q��9?,P;���_f�y�D�٬wj|�ڟ�.��2�������4�s0Ǿ�ڣ�B��_�C�\��q"b.t�9�����՗�{=U���K�C����;c7[w+�1�8��c욨t݄ׯ�/Ape��h�x��`ْ��U¸'��>b0c~>	��!U)��,mːc�"6@��{���>����=�)�r����w�����a������f���>��'�����*kp,�&aè�X���|<s2F}	�>\�iO�� �D��F�ّ�t��΁i3{�������W�.����8�{[4j�gR/s��H�G��a�W>'�i�,��T��V�9!Q���4�Rx(Q\לktR�N�O�M{�^+r��f��~��Q���@��s3X�;�jF��kעE�^"x�yU���otU`�;_���Ui��٫�td����ݠ6�P{���!�X��ߍ|�4�&�(<(�E��+�Qb(�}1�y�gJ����w�̇������������G+	��=Κ�v3�,�!���� OF�����cI@x�2�
'�70�4ѳ�a��^]�K���$�4;�`����a�&��s]X�d�0���7�[vI艚1ܔ�\�r����J�)�+��/��/ngW"e��BQ�x����z��H!����}��F��J����d��y3���PK|f~��	�~������s '���\.ԏ���fN�4W"ƗEٗb��$�D�F^"����<g�>�Ǵq�8�f��T" *D(�����m� ����Ii突�ư,�Z���U��yT�NSJ�;X��#J�|�]/�ܐ��G���ią������_��x>&2�Τ��F�"��1�P5�W�tC9˾Y/�v�dυv�H>���Y���UrP���&@D����Ҹ��	L1T�;,��N�%��@,�i`��.0֌BQ��ũ)��+�8�;�U�i���۶
d�y�oyE�v$G���6�c}�	)8'��oS֌݀�vb^`�K��R��N�� ]��wc�v������D�*9Qr��zt�D,Z��?���a���:�<Z(O���U6�l�}s`�^rw�ME\��ݣ���})p�"rձD�$��w�c���M[v�~c�����=LCL�q�@�� �s{Ov��e�/^ �p���mu.����,�E�0�F��0۟��XT�2x�K�:�l*�:5�+����'ii�8{d8��X�Wi�|3:�>���V�GN߁BA@G�q�$+���+CM������<��L�����E `�4n������:nz��� ^i(P0��aZDq�#��($_��_h�M+��_|떼�r�<��>���bddk���T��s��h�)�F���}�Q[�"�?�Q۫�n�����^j;�ఐ���Ϛ#@�5͜���[��KS5q�� ������78���HF7��2K[���ۈ�<�9Oo�X��+��w��Ɯ�����:�竚�=���i�dX� IQ�w;�E�f_i��S�o���@4A�b��#ε���b���C5;���X�>xx�\�n��O��tc���;���,V{Q���� �ef�������Y��xE&T��z%�Vԯo�u'݉�)+��k�6��N)u�籵��#|tk}��0�?���l�դ�������5y=��`I߫<%���Q�E�
5��9.�9�"w�.8O^O�[���,ؗ�5���Ψ�O��yсʛ����UN(C��t+yǷ�ج�+XT��}v��Dҷ�Kc�:X=4U���w�a�#0���Z����κU��Hp9����)RgQ�?OC�y�\N'��HiU�h&�P�_��2(������<Dp���|�ᚗ���7�1��(�N�:ep��d)a�����!��u}�*P�j��r�]�{�	j�m&u3�f��Wg�t�X�6��C�8�m���䀲S���?z��é� �xϨ�rx�G>��[x�ь��I��준K���2F����+�Y���pϩ �A��k�����?�X n�9W�<�kF���N2���v�e4��%X�������mu�"d ^J��R�o���o�3��6��8��oc�o��oWh?y]|�8����9uo4ґ-���������_`ǱɆ�^v�i�EJ��)T���%�{܉[�vQ��]��a�"���(hBB��|QI�������E��Y#4jP���n�~q���W�W�Z�*=��U*�Ѡv��RԺ��_+��W4�_�k�����ΨW�u����B%���� @�tW�V,�>���
���>���ͭ�i^n�X��i��V��v�k	�Λ5���x:�i�&��ƿ���giL7�7dꉐ��Xn�?`�!f^�˓�d�r-6N�vIq�R��|E�VA�oy�qPf��#$�=��z
Y{��Pɞ>��ۧjU�����ԑ������ҺX�+.�xTVpU��Je�;�e��('h��$����$��{W�	i����$�^�!�'������f���������@��I���]Y��iB��J����s��u������ނ�X���ÃO�V(m�ߟ���).�8X�	 ��"P�g��cu�fq7��v��˓x_��j��r

��8��x�d�+'څ���]ă��n�~���B��r��w�J�S���l����ń;eڭ���2��|�8�,��+\���B��� a��0�+oXK$9f6����P�\`���P��s,?�P�1_8��c�0%��b�t�$]�)
SFR��e�#XÜ*r9�p"-�.��~��8"�k�M�C��C�_��l��R���?�F���	�ET��}~� ���'-vN����ToF��_Ȁz$��ι̯a.���,ހA	��`	�M�&GÈe�C��\�%�f��6q��,��T��B-X�Eڣ�p�m�?�	k��.�/L2r6#�����{7�b�(3��T�d�H-0��UF�:2/n��"C�*�~���XC��w���ܥ�����fy��a����Rlp��5�)׌&$5�)v.Τ��].Oy�A+���p��������(��v�L^t��d��uc{+Q[��#F�����Ś�л�� �+R��L���K	CY�	�cyXO��O��q��
j��K�+�2E� )t�]�5�bu��2���8��OGh����7���������n��uXT�����*u����νk#K��z�&~κu��6f��@}�e�)�k�t;��|U�_���Z����K&�6��:!�}�L�P���	�_h���?�PU-�C�QH\^H�
�22�]����w<Ir�?9cf�r��S-�ҍ�%��yk(�{�r��P��q(H�}�Z��Y�~-�W(���lt��P���i.;��G}�o
�g��b��:���A����*���o������|#���(D�x������8"����B��=�e��XĶO���Lj��5�Z?=c���=���3���-ԋH�	���Cx�k]�AbA�����^�_x_\�}�%�o���86��w�fxܰ������g��뼠%���Vůx�
��Ǫ�'_m���U&o�A�����]G}"���X-{-�}���"�4�}2�9�U�������^j��FϨ���S=pY��k|ҤB��#�g(�wlxjvd/��V(?x��	���(X�$<:BL���g��0>�xUhsŷ]��$z�h폡3��b��z�X�3��a&1���X�eV㕦͎�w�L9fS��_���F�
��-����q�r�GK5�)V�<���g7*0�l�W^E`���[�$Ӓ �\fYp�k[�-i.0wj@�?r{#�\c�h��ؓ(^�Q��Xa�k���)0�ydDy��JqT�F��o��>r㢃S^�Vl��Q1������>��M�C�Ԯ�#��7�_�����F�
SsZ��ˉ:Z�x�9	Z�QT��8�!TK�8�q�vK�(�r�E��	�>L�Dx��:��ΜG�{��4��X�Xu;	'��%ϓ� |�۟V�:��O�I��J�y���Z�v*aIe���=s{ן���~"M2���]F��/�������t�Ƴua���f�`��|JB࿡2�8Tb��@�Q4M�gw��9�ػZM}��l�7��4J�۳}���=��5b%B�k	��<o�UI�d�V�C�\��HoFZ�1O�N�\+���
�졊����Rm�EB��a����;���ˋ��`@���e��P��Q�v y��L
��dz6�K�CSX|_W1lLQ��`m `2!%�Y{*@�RD�V1���Uc�ljom���i�p@�[���r������Y��$����+���s��+�^��r�_�ĩ17���\M�e�1U�l��j% },���կ�+�8�MXS��XL�"�a�BA@��7[u�&�!k���h��s�_�Y� �m�
jb(&���]\P�ȩ;�4J��^��w��vRz��:P:��?�\c�A�`���}�milC��1m��+.3!5Ė���{��<Q�����u��Gm؎�j������go<KH�o�B>��9�G0�(���+F��mO���*
�.�2(}pO��5�R��8+�~���@N@���~&�����B���}���d�X��.۽,+�����^6ڿ�#ܻ�L���������Hi��p����3�g����q���P�t�)�h�Dͼ�P������VY��X�؝[8W�@ ���(����~�·�7����?��n���?��4�D+�?^X]5`�qr�*��r��l��ntתoO1_e	���&0O(�E���O���;�o�[>t��$6��ҰXG�XGt�WF��Ҷ���۝x����Tg�g�?�83����6>7�Z�>|��(K(F,�oBO��aH�v��+Z��Y�/5���A�x���#-�6�#o��y�	,�h�u����@KvONǵ��O�-��/%��������[��7%:�Gz��6CY��Bz���D?�|Ŋt��[�����X�JG���:�Y����C���h��,g*�$(Yx�ze�\�!̄�Ll���L���C�@�����tN.�P����o���[�S��Zr��Zn�:'���h���d��8�����S�������N��
s�O��-��0����s���EgG�m|�e5�Uʲ��[0�
�Rt�vm�W�ډ��<es#�=�4���[L����j��J�i$�G,�L��*�L�(8=��gȽ��.W%�v�U��2^ �}^�����b�E��Z�+፱ȋ�J9zv(�%=�������T0k�pN��6�Z��+�ϛ���=�|��*:�
����d$��e�GA�-�~��8�!���UmW��^_3}�Y;kk�8�բϚQ+��� �R��!Y��q��v�)���[� ��s��m�9�W�������J^�z76�*mZ�;��;��F�).0(o{�*�յ�yߠ��I���G|������3����� ����{��C����W�ٚ�V�B��И��Y(F,8[|�f�~�q�뙄tG1Åĸi�+�(E��1������o@�d���#�Qx`z�t;KM7⪳��<�2���w�
�M�J�v�)H���y����n���4�A�h���1�Y������돢���2U3� �]6��`�O�ӴE3��K��G��eئ/��a鵠d��L�
�P��4|o�N{�D1���D�{���;����I��/��)�o�%Y?$� [�EJ�$�������U�j\�:�%>��o�?���g�:kQ�>߷z%��0�>&Q�᯴�.=�����I$GgfC<�[ڱ}6�r�4S�����>O;�&�v
��j���<����lf"�d_�y��ñQ��"�jZ�A����	¼�+-T�M��e�}c	Q��d��!rv�-J��0̕��NãIMZmrt�3E˶� uNVbɞ� ��ْu�R���/;.���h&ڇ=
�1��4���V>w�e��˦��Se���*��"L~	�_�K�%*����S��k={�5 ��Вt��'��\��e�z�Ս�/��3(��Itx���D�Ҹwg2G%�Du-"d��Մv/'E��Ǿ&W�<�Zt��9��c��7,ncq"�
�
s���y�,L��� �J"�=u�����VHM�آ祅(/%PxD�����Od���-��������u�����U�k~V�p�'e3&���+�U�dv��Q�kN|�f�G��u�g�x�Ԇ^���X��o��"I=��ri[�m�7z��������`���蘕�k�Ú�)"�>r��G���ֹ���.�Hk����@��y4om�E�T&�1�\"$~�֙�T�L�t��p	:�TF�uj7c.��l�O�Hw��.Y��mL�࣒Yx.]�p� �B$�R�����ғ��o~~
I��OJ*/|���N��xBDԷ�[??�U�ϼ��ZC�����c۬R�Y��΂69K��'��W�qN��&�����d�@% ;K�ϥ���\"�ݩ��g����vd�~����&|%gH7$�?_s�{%�ZF�D!H�v��D%�>�0cj\B�2,ť~6��>�|���t��@��d��F�<7�N�k��R,֒�m�g�ɖ1a�*��yT���Y���d~�1�p�=)���1bJ����p���C}[<J�O[fY3�rճ��n2�����U�4^�}��h�R�Cbx���j
F�[���z�8���e�E�r�Γ��@e���)o����ߛ�o�������K����"}P&N�iF�O����I������v~q����a����P�/Aa�ϒ���_:OAI���r����8>��7%%v��oѰJ�ˍp�B��F�ͷK ϝ��ȩ%�-�@b։�7⻮�s��/+�޸�A����,�l&D�x�f��R-��P�9�w�F�P���u�&�(�)u�i���b�Qn���ʬN!�uZ�p�3�����d~�pnt��]��V��6�h#�HtLw�|[S�v]���$vsU�?���-4>,��2��4�R(��'����
P�Z�V��^��j�iHb�{��p��b��kW֟]T �LS��:�� ��^c�PHBĈї�VD�6赒����tJ�Q�O�|�nC���bѷ�(��A=-tˤ��Y�	�'b�L��yOC?�g�*Ţ��8�	r=\m.L�Ky`�Z8����Tb���f-ry�Y���u�+~����,�л^�.X�/k����0�>�#Q��ߓ��˿{��_��nCwVz�'�"�Ugu�������n�Ds���BA���\5���+?.�@�~m_��AǢ��w���U�EgG7�5�ᅺ��4F'��Y��P��nճ�?��X� ���&��;���~��8�(H�Ӎ��˔���I}�R�|ۍR�{��?~�.|Wr
5�~k{bk��$zA�b��}`�W;���wjm�'WA�
��b��&������	���'����wc5D��b�}v��E|�r�0y�����?ʹ�f	���qN	:�l(]�冃ݺ��z� ��q��r����?OҔY�)����_�v�vu�@P��+ 0YR ����K�N`��H�ˆ�!�2�>�C�L�x�&4�K���ݖt!i�%9�ϋ�r;1�������Ka����y�2�1�O��u����;�b���R\�ҳU,�����%E`0���봴���B�}غ/.d�\h����$��Mf�`�W�O��g����7a&|�|�v��Sg+H�C�B�m���d��
<(J�-;p�#�y�dɗ�Q�[�Mpa��L��m,�����JN�E98�e`}n�g�^ף�[b�mf�ct�O/��![��w�%&��}.`7u3&���F])����I�������g+ߛ�)��v[Lޫ��L��Pv��4a��q⪐�L�o��!-�E�!��[����8�1+�44��Z��-U Z���8��65��Hzْ��!�Q8 ����ό�ԏRHb�8/��*���eE�b�[�Z�7?��;B@N��-b�a��zx
��\��5��}|��"NX�Z۝sb�5=��E*��'�ߖb�1Mtk�	=���V5��Y8�A�RL0��W�s�Onf����%���C��T%L>#<j����[G��.���L�џA�4'R����N�S�[i��<QCt܇"���~�8�d�c��y�ɡ=�1��잢�a 7&��R�?*"|�]�����Xp��ۍ�˓W렆��g�RQ0k���W��ɿ[c�)$��[�<�H{�J��Ս(�0��Z�5W�a���{rI���f�!��=�����6_L�i��We�WN����<#����Y_9ʁ׫���H�w�\�Ml�r.�2t��0��τo$@'m� `�< ��еi��U��SI��O�A[b�pkrA��vY*b����D������T���d���+�m^��cb'�i���4w�e{����B1|���俌�&�;�Lo��gB<;�~ROۙ����EyW̝��%�����>A��~�ȧ�Ō��:q��h�zyˌM���Gt��a�ἦJ�.�����DH�7�*�@i7]�U���#�g�j�.Bj��Ӭ�&A�T�7���
�����`:@�J�A]�}��)�r8���쬝�∏����{B�,w�L�x�[n�.�Ȃq�������,,���x���=����ǆ�Ia�z�;Q/�$��&'f���R&E��XRQQp���v�Θ���!E:��+Gy���IK$Ңs��ѡ� 7����^����q��R|{/��%B|[Y�\B� �ݷ� [�Sº����*���OH��Vo�ow*����w��Zg:�{r�v�q^'��?W�(�K��#��Y�@%����Ԣk��>DAC�V]�b��UNW�������4ۨ�r��+Ȣ�hr�X&.���]�Q9����W��vد�4T�Im�>�.�I#{�L������ y!P�����ua�/�L C�{�e���s-�(�,Y�IY}����v�������y����ޮ`\��2�����SC࢕9٪��Ş�k�,�A��|;!�+���f��%!/m|J�J��d��а�?a�2���ƒ�f�{*�G�ee��1}^�|w�w:*J6�g�g~2��x4�$��1'bW�<�� �'��d|�|���+#�r������%5[���e��P�0�Qs���J�L�8����J>�h�P+B2�Q�����l�$?B޼2��D�J$ն�e%�&^��?����� �F�$J��a:����HV]n��vH�y�0)}��-�o��6I�Μ� !*���*܉B�c�j���X,�@�O��nvi�������¯�C�Z���v�� �d���A����ߢ7�о��K~���?���o���Hv�� �k��o�>��0�QQaZ���'O�5;:c��pr�Ԅ�@@�[yg���MG_�1��N/�M��#�����Ze�8�748�>���f�u����B��Y�l�Y>3Ba�c-����P6`�Sf�dth�ܾ�7X�'JHC���G-���~�Q�sa��BV�6:Ԉ�0gʚ���v�לt�!�hgF�-��K���%_rV�kV-eU�i=P�≷��6�R epV�#Ѩ122����>dV�T�x[�=P�"��Yk�q����hv��N�؊�7���ӳl���{>�-�̿�$)��i;�7�������@��y؈�*'m#0m�ï��������H��ٱ,}@�-G�p�u�A��U�j�u���5�T���*b�<d��ꒃ�ӝ/|b{���b�}]
�F��x�R�S12��fI%���H3�O���n|͋v��Z�jMϢ����+�����Mu1�1?՗�Ɓͫ�71�m��`c����SGH�Q��c��=ѦT�㹤����d�!q�x�����[̒���.y�8|Y��_���9֫�3 �ϴ�����/������t�-��o#1~�����"�o��!ૠa��'u�Ƴ^8?> '��\��8�IKX�!9;��4��E8��se�3�ʮ�W�eazgzL>@2EuI�e~$A3���!e�ex�5Ԭ���}YC���2ln�F�荛@PKpx�spᴆ��Pth��_rnx�,V��Z�<����{i潖M�04{Z�ro���&�?�N��r�?*������b!��9����&k��n�1I�	^��$Cv���s5����M��,�k6���͡pX>sw��x��ޞ��95�Nإ�k`�K��c(Q�SCW��OlѠ���(�}m���kA�U�`k����5��!wc;K$?|{��h��\z�a)ؓ�h	�J|���w͝G#k��}�?�o�/��UQ<IJ��!�I^{�o��PQ7��[��(T�3UU��b���84�X�2%����M�mb�������e	>q��%���=5&i�j+�:j�����韑��N��N�����𿔵!�I	�ktN�W��`����^�_#����wU|O��P#HOv�K�g�gXM�I	ݟ?o�˖�����bxt3�};��g�z��}ސ�~�X�f&�U�����mp1�$Gw���Q_Ӥ�h-�'imhH,I���g��#$�\$�1����8	B�\PJ����sebR�L�04�=�_����n�Q_k�h�I�q�9��	�]�Y2ڵ�B&�������,��q��/ߡ�����Z�F/̐�1c��Y�,YTUĽ�������U]Krw������G�<"�Lnoyq1b#����-��� rgi���`���k �����\T���U��9l��=D�lB�%�-�8�-��!�������Yc�=���_W��:$8:���� g;�Ԑӑ��S,@�n���U}�k��wѬ���/���z�z��K���n{2&����:W�Y��]�u2���k�Az�����zEB�4���v]�X m.�%|R�i�9%�P�r�'�*���h����?�ڒD��="*���9Gv����	�㶤'�w��M�5�@�Z/��m�����0�3-����謪�-���r4=���'xБ3|�OL����N�D�s��3}�� MQol�E���)�I��`YR�@�A=a��L"fl�V����N��9q&�I��\QǓyU�jnS��`I?E�%��vk[V��j����e�f�����m�9��F�y/��qNɸ&Yp�X>�7V��%W�!�5��g��v9�w��T��QT�o.Jh������C��{��
�9U3Y��� s��_ʥW��	T�k�f��2S����d�1\������tz��Z�����Y餚��z�w��!)'KzHn<i�3-ً�48 rX����Y�\/Xp� ���
�&�A|Rm�`V:bmuF��h�/)�a���6t� |�n� ��RPh�h��x��ǂ�@�kz�0bܙ�xY�����f�x Փ x�3J|�#/dڛ[���@�~J8��ߞ�sV� a(.�h���ぅ����ZTL�c��[�5ݿ������Ub��
�����դ��Cb���Uݫ^H\�Q�$H�-fd���R��C�?p �,�.��a��!ʸ� �������X_ތ
�M����.�Z?۷�D�����.'2N��\y3�{$�<�����9�Dn�Ε��C9����T\
�l�s��y�i}8�����K�M`�'W�J6X|L�[����t#V��/bF_c�Us1��SbXj���:��o%ʍ�g�����W��'B �L�e�Y�����k�3tW߉���q��W��z�<�7�1�!8_QsO�� L��x6�P �̾�xY�/2� }����U&��F
��N'͹���FƦk�����ڏ��!b�>�����>�(�j�k����_����p&�A�TD� �:А� F���+�#��T�k��PB���+��M�|��&b��o�=r��B�6�^B��$6�Yf���_��<��gܙp��ŊJ>�T�]�%�6���uͶ1Z�-������s��]$G%W�p�+�@��0��R��L"�*&��u�����wdG�" kÝ,�8l��z�3O�CN&6�ߗ����9s_�b��!�-O�`���P1���l-���vb��:�5�I������F�!D<N/�n�"�9>�Ob8��D![fq�!4�� ��wty��H��W�B>�n��@u��t��M����1R��`8���M��M��Ry#�]��S��b�N�Ȋ�d�`{�,ðwX琫qJ��7`xwFJ�kz�A�8�k�?coc:[����Wl�	�����?}8��{_ L$��9�1y�y�r�l��rD�_�u�G�%C(��p+��F���Ғr�nF{w�_�ZF=!�Le B���C��2����j �K��f	(U���g�|.�S	Uf���y�=��VQ��|m����v@n5=�(������8���ʀ����,�YC���_r�ђ�G�O3}�R�+�pL%[x��]�U��]k'H���(t��d�F�g;�aZU�yC�I��+�a}��@@�`�H���؞�v;���`j3���JfH��y��ف`.y=ed:6j�'��/�=Vt�}������]H��;kl�m/��8
�2���|T!HX�ƾ�n�G�R����� \v7ZBg�-�t�X��b3'?�t1�8�U��_L���@�������B��-�w�j<�\�����L�1�4q�b�����Nts�*T��숲C)hPC�D�ix�i��#��5we֟541��^��%U*&4]��|^Q�㓗^��4���S�@��i�{"��G��.��E~�?P����i�ME���Q*�Z��#�և�:\���Ļ`w,�Io �ʏB��=<���T�	��֛/���E���
�I�=B�}*b �-)>�?��N��`b��/����m��ZP���Q8G)�TC"�f��� iw��H�2fxY��&)h'-/�ٹ�{O|���ݚ��L螉'z�-cv��GJ��@�y�ݯ⧀��V���"�iK�������1��̙&�3-����~#s&1��M��!�������l��m칚��1
���`3CaY�����?C�&Ȉ�0���<*DuCK�����+��kц����~}�����U);�ւ5[��6-7��V�5f������rG�~���T�*R_2�-��6'?'�HŒf��@W�������58H�9�D>||�]�7��3$���Z����x����B ����E/�q��شlc� ��Jx���ԞI�7������N1�n�ר)%��@f{�`��5D2�	Cs����w=�$�. Xs"�a�gW�$S�;�ZR%-��57�H��� �VO�Ї|r`֘�/���5�+�cN������x囙A}��W�n�Q��Sg��Gz.-�N�7�;�se������I>sW������7c�/�SP�<%����� ��4�DG�_R��޺�E[L������	�e�n�	����oU%䂇&dK؈n]gy�?g��f�Ƙ���N�6T ��oܢۘ�F���fX�c8s?^	��:s�����L3C<_p|�����J.j��#��7ޞ@��|�|)d0�ܗ�~u�#r�f��p~6j���q��w��n��7��.�X��4�e|Օ8�X�:T�\���.�2 ��`"L�C��;>n�9K?��oH��?jA������8�Rϼc��ϲ���vѯ+,b��c��*�O䔋&���!$����C�9�[�eqJ*�t&$���Q��������_?�h]NV#=o�$U�ӿ��r�=�eX1��'�0+����1��J�΀�*93Z2_@�����M}�?o��J䟑I��	��m���G�� ����B�a�w�)!R)��^�2���ds���R��F�K�B�k�E&�,ϑ�W� � �V�<��OZ�Gui�7��=��u��D�����Ir��"0.�/������w0
�c�ꈿ�@^�S��a��C�ފ�[A��e�zEK��[%*t��uNh�)mq*Q奒T�IB���Nh��֗p@]�е���ظ���҆E�j�ๅ2gba��x�_E#+�8��L _�ɠ���F�rn�j������_@�7�f�0��p��R�hܣ_bU��Ȱ�F����v��{;ku��W	��6b�����;
vd��<r:_>��z����U^> a��;-����,�#���X�j�ܙ���,:p޻����x�	�jp��1��N �_۬Ր����.%l-�
��q���J�.���o�^
�7�ｄ�f�S��plSa��.W�x3��HT7Ӽ9�<8l�Q�j���*b+�ji��w*���,�7�w�J�o
�c�1�}&,a2� J3BvE7~
�Wy>v����}P|��d�Ls�G Ο!}̤󓸀�B&e���o���(��Վ(C�F7���!0�i+6�%�!"�ੌ�2���)��8�+�1ڍ��,���|�1T#� O��=7�Ut���`F_n$>Cb�n{��^Fs>�߯����3�]?�����fB�3��hY�Z��?�m���/��:�`�F�J%�b����槊��"f�2�5���Ҷ��.Q�»�T�e4 J��z�K���>ȯ�K�gK�{�V��v��@T1/o�9��1RF^�Cm���䧷]iBo��3���`��.��xzWe\B�%0��U��ϻ�v��÷-W��}�UY��~�uy��.vW]���8��4����� wVd]9u}���F�@v�h���⏓@�%�<��a8
B��E�~SۓH(�w�F��H�$[W� ��>���Go+�qby�,9]gdZ�Twڲ��jA�����D�|�Ē�V�K_I����N�0��1��Hޙ����sg
���PL�l���UD��I�wJZ����8������vY*��d`�X}x� ��{����=<_&b�5h�L����u��(i�g�����~uM[�S��[��;~'�Ai�����/��n\���Gr9C�X���Ԗ9��R���>אۻs��%�7�Qy�s����јWl��~B�_Ý�,A�xmi^_O�=��L|"V���2��kP��_|�o�^�hĂ��:w�QV�V�{ ��}�3��ڄ��:��/�P�.��9��"���,�aIp&���̅[_Hf�i�Tl��c��a8�%0�eg�X73� 6V�ⵓ�3�/L�H;���aB�Gr@F��.��G�`{h@.���/�h�WY�(�iH�ۓ����"��!ş�b,�s�dj()�L�����/^I-�ұ���. ����;D8h���6�y`�؇�� X����R(��p?7(��i++�]���"��R����:^��-	8�*.N�q|!31�~�ʋ�Inϗ�z�y��[)"�,K~�\��9�X��2���8�ɷ���Ta�swCƖ:��he3DE��exf5�����+���s0�^���s���~\�?�dJ� � i�=/�h�ç>)��5%�~Rʓ�D��X�ؓ�����
0ō�G�F����?m鈷"ಋL��	���'fچ�k���	�p� »�a���@&��u�{]��y$�2hc�_*��+V���C���A�^}ۜ�O��6�4��}��w�s�Cl�Yb ez��g�����V,�c������t�����t��l�����Mʃ�П=�+{Z@�<*���#T��mmH������0n�xX*3�0I�6�M+X�p��Oi oڻs_-�<s�>�q@.��w��`�z���k��ƪ�ޫ� ��E�0|)Cx���ǑDKݪ�:�hUzt>CW�`����/o�Q�c�l>B�ڼ��:��؍�q�7g�I��%�^��}�eC�]EM�E���E#ni�r�rN>FꞞ��I�̦��P�����Ѻ�*p������T��14vߑ�/��������y�R[@��;����{"L�>��jbC� ����{y�?��&(�t�����
37hol���U����(� ��`�&�qN>7�t��9R��T��=~����h�bd���ۙax�����D�<�7y��p�Sӝ��o�W����5�@(���喤l�k���}�����1���1��y����v����xů��
��o��5�OVx�t�4h��s�}���3J�]Ӄ�b��z�L�~�EӠH*�p|�Jp��·��5�/�Q�=��z��c��V_�V"/&�@�{vX-I����ß�[�����K�3u��]�ӂ�+nS�D5~��K#$oot�hE���Qڱ&�'a8�V>�����4�R����T3z��=Ff��=���C҆T�,U�O��� ��!��qEwy��W��^B]�xr�3�ږ���i��k��k�^F���CSjL�c��vYbfP�-nKD[!���~�-���������8��1��t�o��ƔWw�6o�E�&<@�r�g��Y�X���3%�3�ʁ��::�O��M�D�f���yHM���R�J�=�ާ��vtO��D�LFd	�M�MUGU}���d�G/pZ���F`�Wx[�2Jh��E���U�<����IP�Ɣ�3,_�G�D�����T	��p�r8a(��|L�e�S6��ү�4�q�J����j��`��T��~R��Κ]5�y�b,�뗾`�f��ǗtM1ے�����ep�	oe!��p��M&���p�#r�՚=���F咗��z��D�"Y<9f>(���G��x�k��:��n����� ���Q@G��jl�L�SA~��M� 'kRt�(��G��rHc�rWӇ�ӈoR�{�T�A��D��m��.k�������/�}�/������*0�/D[��[�}��T�P�%N��'�M�&��(��hr<.��yD����s�q�5�G�P�cƩ�k�bD��%���tE��	�F�d��?�a֟��Y!}�Ɖ[�I4"�m2&[�D����^,�!1:g��G� KFoO�<-ψV��mj�
E-+�AyER�9�6^��#�	X����-�qe蟮�BȜ'��7�TY��Q-��/�`�%e����^��[v�����;ͯ����W@�!h���"6�v�7�cD����>. �DD4f%Ӫ� �X����M?�s.��9�b=x��^�'H޻�w%ZT[x��+�\���3K/���(_�a�	���L��[�
����Pa�8f�p�ί�o���v���I�i꽣TH����Ú�6�0��Jb�W����Zf�]�Ϧ�`#�õ��j�O���O<v����sύ�*q�v��{�LR��<����Y`3�\Y�\���/� KP�+�֓f���{Zr���"�jJ��u�^TQ�ۤaMʓ����ؤ[�m���+ZcU�8ȧ�Ay���^��x�yN�HD��5߭� Q~��,����"���.�s���#d;[}GE��$���L?]|D�^�>v���8lf��T6\`iY��
�VB�}���/J�����XRg 	��z��:w�����wcB�����e��vŔ��ĥ�:`|��w�կ��Nn�r'
R����` �w[��-Z+���i����/ �� �s!�� d���:l�ZM5�C��V$���q 9��Le�<�@`�@7���`	��s��ߗ�0N����$��q�L�>\I�sjĿ�D�x�_����/qȁ̏�S��;��K�����j/9��U����Y|@��zؽ�q+���9�bi�J`b')�����_'�DB�Q��cm`^*X�g�"9ns�x�k۾��l�.����´Ψ�$�oBRΗZcv�C���}��Q
N��M[��� �N	Y���rF��U��oo�߃��-��Ӛ\5g�<��-V���3b�q�	&�I��+4�3#0���FH�1J�F��O���W�Rd��Wr�cw������L�Y+��;����4p�kF�cs3�G�2:��)6^�R�H�G�|xc�Д��fA���<RN�\��v��G���A+��Fk,b�q��n>�*c���8�VE&���.C-�ǔ3׬*�C��B��e4_D��s=vѮ��±�k�!b\9��Q���15u�G�:u�y���^�����q|w�(NoʈQ&�_�IׅgRč�ԲI$m�pr�2u� �K�UK��F�6�P�8��j�"\�
�&;UW�,�d�+;B ��Q������z��\��e�@m9�*���L����n��ֈ����bG����K1;�<����R5�B�K��_f�������XI���H_O��2&�>�
�NB��By���TK����	��i�Ì��!-}��)��/d��,޻?�d��C�����j��ho]K2̉z��R�I��#�D��+$���c���զ[tןӿ��Z�������P0M<9�oD�_]zyf�9fD�x��Wb�~��s�MF��?z��Q+r[ۤu��P���1��k`� ��n��Y>��-{��|A���������G2Z6��x
4g�w���
g	Df��y�����M1�8Vw��<v�F�m�8����Ư�Q�ιԕBЀll��{���'�#E��z�T��`/0������;?�`��a������遷e�V�Z�̰ksl��:]FV�m��(00��?$]����Aay���R��}S�}ܚ��V���+�u�<�c}z_>F���>/�(H? ?����R }�o�vUm�wk衃�������{H4�~=���I�f�@�}0���z_in��CiH��Y�B��g-��ٯ�xW��*�od�I�����I��1���)w0y XC��a���U;�
�zJD�24�&ڣV#�~����F��[����N��ܰMhA���3���֒+h���R�m\��{Su��n<zR���Y�Gk�J�|�b��uLoxB(����|��Q�bbY$��У:G+^���֪A�(��-�Xvx�w^m�T��)W�ٯV,-�_���-�I?�Tw���6L���G~�៕e:O���n=W�K�^�����P��Ы-����-�"�ڐ�$*��̨��]Sp�2�k�D��'�؞�������3��O 1#�9�c��蹄������`�ß2E�m:A�ƯΒ���+��^����� FeP�J�i�Z/���
�SsB�
)K>2���,d<��QႤN��I�k�,���I�A�����]B�JOJ�pA��}r�&��6;D�M�V�	p}� �i䪵-xW��%�����zޕ�t�6W����0^M�6m�>g<���ޒ����1�;��e����b�S2�1�P�m@7��5d��\�,ͨ�yfX���h٭�A���h����dE7�f�CR�b�Q��<��;b5��4��قae��쬡I�n���f;_|p���ڰ:iѰ��y������MG�m�j�R��`�4K��$N#�+VKo�m��nt�!��B���D8�Λ�����c�`UA�T�M�Sfn-Gв�4�Q��n�>�a��G M7s�e��aʌ�19R���{?�46�M��ی��Sە��L3���P�k�=���,%�z��3$�!b=۴5(��A�9ݹژ|�M\0KϺ��<�Y.=�br.]4�b�t��)��\���pef���ďuP]�e�0?],rf�/^ݿk���XB]~�I�D���?T���`dk�!�]]x!J)�Nx�;���SnB�,����(?D�3����&*�5���@�|A~�I���� ȷRi1]�$P�W����eZ�����~�)�ɶL�$��+(�Y��=��,*9o�ѵ�Rz�bQ���۸�G���_5��w~����I��r���7!�9�>Y;61��F����{��=��W�,V���@���*jj��=7��3���^/�=m%PI������O޵��$�7|zw�?QE(���Ų� �~�慣^܁A�QTp�q(g�!<v�L� �,�����O��OQ���^���C�����5�9�@bf�C#��~��v����'���X�;�n<�z�Q�G-Q�piӘH�MS\VY�M�͉~��D��4>�3R0[�k�3!�$��It���r�/$P?�?�B��s�O�)}��U��F�E�����z��#o����\�쓁2�C_6(��%�Np����e���ya?5D���R�D��B'�����¤ۨg����u��m�r>�8��#��s�-߉!�IJ �: �nAQ�^y��Rn���<���w�F3"�64T�߰ʸz~TF�����nW��wx�G���:�䪎�
��>�I�o��c{�3�e��,*�C��_�Y۲�d��e1x�k=���ԙA9ҏW�n0���ض~�Ҁt�@��h��Ǘy1�y����c}q��6k�m�\}pǖcf�5:������޺ϙ�ߛ���qfP���ǏR-�������R�
�Bdvf���;��1M�I�^mW����>I�t��s���o��\1yOW/�?`H~RI�o{�c���& ��) �k�e�����*�D8�1��8�\�����w�_o���H�Z{\��l�@P��w��M�W��� O�ӏYӆ��l�@<��Iȩ�w䫽څ?H&�j
*U,�`�?]���T�O���1j���x!��u>��
�4�Z��E{��# ��;'RT�*T-�*��:KPM3�[Цl%Մq��Ϲ9b�?o>ᜱ!�~�!а '�bWa�Z��s��&B�c�M�M����ɩ*��)h�ҙ5���h����í��h�k`b��=�f��/.?����xJM=X�\?�٢��i����Z �'�/�"�퀷�˓<�Dr�q�T����$ε�p����h�����̎�h�Ʊv�s]as�<ք����1��ylFaĘ̵�{�)�����FM�k��a��h�ȱ�=M��7�+Z�b�>	�q��v(xa�Q�.���~Yѷ�r���<�~���A���~Hʶ����)<���" �Wǎ�E,�z+��,�џ4��
b��v�����/;y�5�=����Oo/="X�fHisf���B�2���.�
Ԅw}e4�Z�loi9���}l�3�nQy�S�9c�X��ܨ���G�\��yɚW3�$���{�"6N���"X,=�
��9w?d=�n����:+��a�J����Y
��K�5߻xz��dV�p�揠4��k�/��d7w��A�M����:���JM+�������A�6ӳ���1�a;����S�}��d!~
*�ⱒW�/��'��r����|ED"��Aʞ �J���w�L�D�:'��腇�H� h1�<���- �؊C�K:F�h�6�|K�卥��s�q�B��qr2(�_���B@`Z3�ž�p�wP�-�9~�_0���أ,�y����� %��mR�
@x(<�N�+�����!�k��Ch�t�� ������YM�s�t6��rY�� �>��f���Å���vٝ�����oضʕl������ז5��H�~-;
���� '��q�R`o�)�Ɲ��y�%w�]|�9�²\*l`[P�*���sj�	�\A�xZ��1AH�L��v����;�D�t�� ��V�x��a�ԁ$����˄Y@yL��F��Z� ���p�QF�j���$�����ð.*:��?���k.h�XB�?9@�R�~���@U�m<���I$���6x["��������X/�����{��#��](H�0�L��E�Z�(�>P�ۏ�"y����ƍh	�4�̆��y�P>��)Ǯ�b�]&�j`��jY��ݫ���7�j�d���`ʲ9L
�,�x ��4s�>|�\���KlE�4�]�C[z7/�ב"��!���0������1_�m��;ޅ�	I��x׿��J[��@A��9&+>���MfC7I��+��&>d��p�$�X���}<c�V�[[h_���L�!b�	y߆�eg<�?."�k�\�ׂ�s����(p���Q�wT�Ӊ!ۥK�wBg�h�Z�q퉓'��R�=rJ2�j�z�0Y$�I�3y�)C���3#A��%� ��+�'�r�Z+F�(Y8�G�^���k/��,�P��Փ��Sy��nb�l�Hns̼�	/9^���2�s>��j��/T�b����U �yλ��q� _�Vu6T4�8�N ��7�%*�xSJ�������jF�y�&��̢Le���/�!`M�cp�0���#릱\�X���Ĳ�?�e�F��s[t�N��͚�v���+��OkX=������ȼ$^��<8|d�^���&�R�����2"ń���b���]�wj�����ک���t���n�\��/� �ɦ��JA���Nw��6ˣ�� ��]!���2�,`�0�V��5Mb��è�%,�wx=S�<���8#do��k=�e�N[e��z��Rɘ�`��l��fWͬ�E*�Pb��C�/��ȄsR� ���Қ�s�ī��������Y���N"}��T��;����2�Y�<�A�eٽ���_�`�#WCCf���4�x^!�*���M)�d?�S`�L>��@��:�����Rt͛f�v{:%�����W��ƘCrSgi�+���2� ڳ�3��褈F��cBNo������ۤ+�T H�+|؀Ob�4��+S&� v�\t s������p�U������2%3Nx`y�\\X��y�"���믹��)���>�`5�*�wXC�}��crD�zx�������=|D�& ���}x�M(3�o���^0��#���SyA`CWDFN*x�}h�I���WM��R:Y����:u�>l���2�u\mu���s���DaX4q�ނ���w��¯�BC�)nZWt�#y��
���p�?�>Y��'w��+$��yd�#�����Z�,����_`Q�5&�Q����T�{� ]{&�����8��}���=�sMZKX3�vW�Pu����l�he�P��N�j���p�}������i�I��@`��;��]�H��_n��,r[,�J���6 �O���3T&l� �w�n�����j�+S���ݳ��0����\(l ܜR8_[������3��^���zr�;$� ��b7(�qI�o�hk�R�1hZ��#�[7!�����k�V�lS�|.��pY(��:~O�f���6\�ӕS��+�/����\�]kq�e�Tpg��-e�����J��C�fB�ִ ��������Qt�c�@�F�@���oͤh �5��i
�����L��J�\+�(�ܧ����"� FZ�֋x�{�#�?�
4| \T�[�Y�?���Μ@���Ӄξi��� �u۶@��5�,^է=�Nv����^l�vѿ�g&�g��Ao�ZZ�Y�!�h=�L�Z����۳R�l�j ��P| �s�]��-><"!5��@��[ԈI�/P�����:����H�fԪ��(�����t֖aN���a���~����v$��k�i"Ո�f�Jҋ�Ù�L�$K�ZӨ��Ǒ')��ʃ9Wu��J#��'�<�YÍ���bwPߤ�YC�̿�-���ɽ$��` �!��e9�b���cF�22_�5�,wQ�rp�_�&�Sam�!�hKÎ�v���z�/�&��Rl��Ta-sB�5��i-�yHyp�Jw���9�~K�	U�H�^��v���O��,���O��@ܰ��㫇*>c@	�.JY���%Y�H ����^�y=G`���>�䟊s���">�Fb�Tw�l��Ō����=B�
���^S�~(���,���,	��B$bp��_R�ih�?�T�nYʈ�%5���ϧV7��_$)���Ob�ftXp����+f�D�Q&�X���Z�ٓ�X����f?m)M׼�"q�s�&��~�X��2fu� b����JA�	���_�&�|ԃ[ g>پ��w�2�;ʰ!��<���ν���|j�{!��K�=Q�����Kb�zk����1��s�Q�պ~��e�s����<�^,\N$���}����#���S�Z��A ����uGP���/5�Mi�p��YJ��gE�9�{���Ut�m뻹�g�|"�冦��q�b�k��V�qT��4��U���{�3���_f�3����2��rvj�4��W�ҕ|��vH�ÑP�VȄ�:�S|x�<�i��7kM�gE{c�L;�j�M�4�/"{��1�=8����YBp}���^�E=a�p^�*�� �]���m�֠�n�K����� v~ۄ�Ie�a�Vbj�&C=)�yo����d�+�7�6i��z�VXDڍl�:���¿�ts�Ɠ�f�k��J�q��'��/f4E�R�rAhn�T0;�"��1��b@��炵��a�V���6����e�ZrnUv[8᧍����Z�Դ�4������f)��@y�ӌ?���G"aF��1�P-��B����*��-�?1u�h������P�_�5�`��`�_�G��`��@�N2c���ڲS���^aTw(��a��������#5�ZNJ#�/dzM����i�J�	���Y��^T�_AJ�b��r4�㘽3�����T�_�������o�zq�g����VIb^k;�9�}s�j��[�i�%�y��)����q�G牮���Z�]�S��� ��:'��E��+.K��8�C��Gn`W�X�-�Q��ɨ:���~��^�'*]���6���Ƴ�����������@����D�2�,J��}�n�/�7#@����n<-=�]��d�Q���D�:]"t������ߨ�����i��7�,_R���f�2 %�"b�ĕP��ʆ��8��f��`R���H:��N��@�@t֕h��{�\�eؽ�j#n2�uҎޓ�).}_�Z�;
�P&X�{�-kn��9�jh��g���|M9��������?uIzubAΏ��P1�1�i��ү�i/�{Rz1fƈ!�ؐʱ3���l@.|>3 ��oX�*	�փ��f~�ai��-" �CGxc�]r�e#��,I��ɔ;93F�
��}2k�����Ъ���X����Ru��u�d��V�UAKB!BA��^�7�A�$3*�)�;:�4���5�V�E-T�'3x��:�t\���8c=Z��?�<1:.�I�&���S�χ��yn, �"�qpi!ND�<)�j&�ɫ�=���5��{-o�G�J�Ӈ+��m�M����'�(��������t��hIv�IϦ-�uA9��'̤�{zV�>�*g�.Z��?��'���� 3��]KF��a�'d������J��1�V#`<ÕYR���k7[0�,�*�F�zc	�5�5�+���wl��_�tD��q�mHמ.ӑ�ѡ�
KS��h(�����b��?�+������<r�KY)��֕����2#��$hAt���^�R:�B	�η�65�U��H�p�Ν[��9�{z�����֔Ka-�ڔZ�&!~^��r�i%7zҊ;��%��;}��f�b��*[v�¬=�72{2���yqE�y����T���Mۡ[m�jxq5�����,��E!/�5%�������ˉ:�d�> c���m��b�w
������,�]�oF0���!m�e���?����ͦ��F��!���\�4+mg���S���,dѼX�mHi��f"�Џ:���>��f�����	�uN7!�0����_��Q����/-��(���Ǹ34��!n��H���N�K;�����sl�!l�������d =��nC�}o�Wf�<Y��x<��dB���7M1B�r��3��(�{��P��8(�V��=}+�-���}�z��!	��C<��4�-���N���?��VjL��S^g�aŬ����oM��4ko_�>����.��S_�����GU�=ㄻ���D;*(U����c"I�&2u|T=�3`�a7H�Vpn�it���(? ��I�ހ�������y�$�%+Ֆ�j�Ա�jǹ�x��f����#B��bi.��_��=��fÉ�l縄сQ�r��/�����1�x�߬��"�k��'򂅑��U���t�Ì�������(�"Y�j\ll��s�7`:&5P�[f�%�R~�a�?~�j��YXG�����%ϔ�Nms�Wk�,K�.�=�v�+�X)�͂������6�9��{DnL�Ȉ�°]'���0u�4S:h�/*p5u��e������(sj�.��`ו&?X�����F�ֱ��$��Ʋ�&��b�6�S�Â�S��?ػ>��k�X9?�#�o�A9)���'��%���I��dѿ�l ��Q��Q�X܃��q��o""+���U��9ݥ���l�8�����8L /x����і�)Q��q	�<�zQ��� �1hSzћ��W��,�/s�/w�62Q�kf�u���L��G#�p/�:�Tr�@�v�( �7�pD*$�W5�	Q�Oq.���	ʌ�k�wY���γɧ[�9W�"4��'K�BVd��9� n8�P� �#[�e��)@:��F}G�U��)7o�K`�}���$:�[,�>Q4�o�9��ݟ>wۆ0��~-������ǻq>�Z=���Cߝ��q�MY���g�Lu��s��XuǱ�~��|��!��(���ֆ��f�#�hC��w�C�����(��/+"��ԟ����³x ���B,d!<��w0i�Ψ�8le!O�|&�R4-�Tx\E?CCnTr�>]��u�ϟ�}J_�z��R�>���?�Tm,�W��D���V�	!�q��d^�;*]���*C�L�����8DK�ݒ��noُ�ߌ7ۺM� Xp�|���h&�J���Ԙ%�Z���4�A��0�\eA��KV�ðI*�t���(=<����pω��g�Rt�VR�yY�?c���n.�||�;�������Y�����{��i7Rj��{;ܲvdJ�Xw�  ��eļ89�b���6Fg`�����Z�(kG�w&�P��&R�I��;7�G*.��~��Z�V�@w��h.@h.�ï�.��\�0Ys�%���Cv9C6�ʮ/�2�n��l����6�\�	��I��6ۤ�{�<�n35��}!Pa�&� �6C�z�����t�+��*��|5��Ď��.A�8��X9b�(^���F\G�Y����,E�v���w�:�7A˓mI(��GR�<�?����f�M�*�΀M*6��k� �j/���c��C�x�L(��<�UT�v%�8��I��[BHRץO��ϧ i�%��˒��p��$�\��c+�F�FƫEk+�I�c���Ə�gMr������Y
�*��|�	�6�/��#Nˁ�n��7��2n������ԏ�:i�>�>o�s]u�bO�ف������s�bKc��l����t�i,�QxAL�r\���5Y	�����[�5��.oN��>��f���İcT]�kԞ�m#��$a/�4��є"^X���Χ�i�����=����,ǋ�lN�ڇ?.�h��!Yi� 1��[�"�W%��Z��q���8q�]�_ɥ�1����>��I��VqN6���Ma~=����<�Y��XJQ;^<�E ��NMܻu\���6眤=�.�H� )Vz�'k��rJV0o����ݧ��t02H4�H|�	���$�������h�=ݍ����S�W͆j^E��A��Zj�\������7&R:�*�Q�.�0��hxx?�q����5r�lƷI�K��+�C���J�l4�4�}Cࠬ֠�I�'��Ka�Zv#F"�_4�1�n4�3Wr����n�/W+�%R}���ژ*�b �}7���"�]��+ �)�3_
���B=x���C��&0-�[v�������d�4?Z�i��;�/���K�Zp2�~y~�)ڴ���-a[;�B= N�? P)��c[�P��t	�>@�lV��}��
�1T`�Y�X���c�`Z��m�����Wz������ �!���Z�XF=��y�n�s�F4��*�.��fZy�(34mT?g/��u�h��&>�[UY����{Gў�GJ'�K�6�z���J �����y���2Dt�kh���YF�o����
h��CyǸ��ugE�\o�i%��.|/��[]:�����K/���ǝ͘eV=^7�C���r�R���JI��@biz�B4�O�(��hؙnV���kӂI��*Ŧ���F�Y�|��wOCPl���g'_��T`N�#$���_$EL\F�\���6�Ԣ�~��GFQ���d��٨ �.uZ?�1����^P�*��]SE�_��Zs|�|ͫ�$�F�*�<?�dd��&�3��,-��(͞q�U>�(�����=���ƶ� k����^!N�_��C��5qXZK
T�h��U�4���~������UW�A��(��	����ad��&��-Պ�އ=ɨ'�V��{����*\ C?fR�=�3��N��y��G��v�i�J�*b�B�3%@"���t��\/�}��1��Rca��Ԯ6�(>PAB;z���M�(�$U�I�8�r4�<�F�˔��Hb��R�����A� �ab��� ��ۃ%rk7]���tX_̍�X�v�4e_l���!>
W�a�7�U
�Ǯ�o�{������}�2��ZC"����_��hV��]^I�=�r���s4g�դ�=�V��홌Q�g��Ps��{��A���^�h�>�/�[��i�:9pF���O�-(dxc����ْFX���� �\.:�uN��sU���~��_��N��t�ˋ�ߌ��t��Y�|��:�y���t4!�%N�y�Y]g�9��CpH�����v��;&Q70u-(CU	`Q�=<��UA�^�A�hR��Ļ�Us-�&�0A(��N� ���L�s��F-��^�<|t�k���e!4�R��8�ꍧ�t��%Pϒ�/��Y_rĶCGw,BL_)~��8�W�I��Q�v�R�G~�cVG2�s���_c�+U�͟T�^���h�z�b��d���cy��ݤ|0����r�&���L���Wԫd�ă�v�����zj�@�N�G4=�S�K=�z`Խ{X�b�5[�h�>�#y����a�B����{�~ij��~����)}��UB��M��3���"�����ׯ�ouQG&�{E�a*K�A���0*��_�_|6��O�-��|�A�5�u�2�~�$	5����t	��%_�|
�o��q������^�,q��9�В��R�_
?P�Λ�)q<6�O(��y�sG������7m���}����Ȍ9��(P_�!��Cl��զ-&��O��D*�-!��� |~k���� ݁�K��st�v��<L9��
�]�$۩Q�k�l�-�9��xfٺ��WX!~����{�o֑��hS�ɞ$��d�����o@�7N4ڲ����
m�a� ��8�.;�	��N�:�8�%R�n ]o��ו�o][ay������e��0��R�ܚ�F���I�O��m�U�p�8������CXn�nZ�Y*�AE�*�%U���>�uJ��=�����8Lr��zE�O�[�%�]C��_�8��
�D���z�� 5y+��?=��\��"����J�Z�d��gH���cl��v탬���s�k�0��!00����ipzS�Ĳ*H�z�3�B��Jȗ�M�J`�.dc�^���..^:�����*Ɣ��!%�nd}�d�l�,���,Ob M͙�I���c�m�~q0���a�荾��ƄGS��
�m;4�
K7�T�-2ԥI���@�Q���B+�0�;e4R��%:iC��0m_��l1Sߵ�ػr,�e�?ɠ��ʟR��������Q�
y�l׷m�B*^�<��¬:]�.��^a����5s� ��`��t����_M�{�ُ�$�->��~�çk���O9�������)�&�@��G5.B4��� y.���n���+�n��cu�G�	���ޑtH!>��z&EG�MO*�sWg�&���=<��^�j�JtG�����&V��u���Y�/$ g��X53|GB;����h�-˷����8�g�?rWyU�`�K'�l!���{��Ќ����8�oC&	m�v��L��[H;q$���I���l�-w��4��_��vR|�7 �W��s@fHɈ\�(�d>��P<q��gҿDCx�����h����!a!��v�z�*[x��5�[3o�3����B�Mf���p�]!�:ҽ�Vz��8���Z�NJ�'H����쀑�С	zC�����sɬ�L����czi��M���(��,��Q�@	+'F�(n|{�V�Oᕪ첓�#�u-��LaڟoA�u��|84�|q����ñ��ۙ"����gE�)ɆOd3 P�"4��L��*��T-黼��c�&0�ǚɵFV� kC��꽡!�M$K5B������?��C��|�?����N� �:�zV��~E��Fσxl䶗�E��*�P�%���=�6^Kê��Ѕ�����#o���_����<J�%�x��(�'��ZKr�����k�}7�}3�ctk��m'G̮S?�`z@��C�R>Q�<�Jw"�%^¶(���4�{�9;v��.IZ[���er��#yl�Y��J�D-b��v��F+x�e�]#����O���`@�+��3)��K�g]vn���'��q-��i��2J�*�K��[�͠��W�Liif�+��z��W^O>�/Y�al(�k�BF����q 4����ʞv�rl�Zx�^�`���5�l�E��5\��6B������N��"���zKkS�Py�ަ&����)�r�M-�.��Ee����P	�D]R�L��"��r�����L�C���9�F�^����mJ����ր#�/&�An�������k+��I��4�9������Q���p+�V����j�����JoL�+�mz��=D�R����z;�bZ�`#��/�B�㿢��?�]��M_$�~���7�E
.�x�3
y������	Z��j3��\aj,]cq��^g�5�%z��wOG�iJ��[�����=v���S2�\YM#50EAzS���ҽ0F���}�Eޘ
�*�Y�*z�+�l���"���2ݵ�����^+�5���Y��x��~|���n7꩷{��?�>7�M���?�����I���O��]л�I�[lfj��x�Ys���	��(`-ٟ�-g^��c'�hY��~l�x����%�#Fe6��Z�����Ɵ����K�Ό��I�Ə� ��$�	g}��Q������kD����E�<I��E�v&�1J'�h>�
�(Z���6s����#\>[l�F��w��#��KI�o%��x�M�XD�Ƕ/�m*>/VQ-\;9"�/ȵS6��R
Qo�8��J#Y 6[ːU��ش��D�p�����a ��iT�/�J8���ɋm;���kҼ�9^�J4��\��S��H��������'[K����bj\�Օ����G��C8`�:l�����J���ţ�#�~�����yV��+���(j�G��VhR-˜g#��?�Kф�b�i���Ð&�1`!����uP���f\ѝ�ל�Y����zf7ĳ8$���M�y���]<J~Ư��B@�O�%E�$�ג��$��55��g�凔Z��F�}�{^�0�vDPXRL0?Ye�μ��R���*��BQ��}"{�t'	����_��xQ�I~�r;�e�P'P}f�>bj���UV�h�-��\�**Y��`�>��nY᝘��!1���[�n�"�1H�RAu��޻{^#ƹ���Y��-0�i��uTa�݆�2��0�^Pt��ː����ŭiؑ�,��N��@~Ӹqg�uHucN~�ֻ���t�f�7�����&�����0�� �|{��L����n'�Ȫ�+&B�]z��j'�Pq@�����&|A
�W�&���������M0`b ��xgf��1U����I6��8�\� y��o�x���P��q��(���? �A��Rv�����R n�>O	��'	�x�.7B��ɾ(��=�3�4����
�������ըZrC�m_����c�{F�#���$!���M�o '��Y"�
�=�B;�u�8�i��34�D����0+�'u���nZ-S*):�Τ&�5����|�v����	Ǘ�WC���ܨ��M��:)<8��r�2���>�(j�V��@L�^�ߞ���%[����M�@pÂ<G)��YL�}V�
���[����r�u����-�7��q��L_��x����L�p��҇�f萎�4"���|��_� �l|��0|c�X����i���-��6�tи�j�?�q����l`���ɟ��38�ФsiN��R��3N��Oj���V�M�A� 3��d��,_	�+��a����lނź7C���;H�ND�T�����oB��;;�6k�����ʅ�E�����g[G@�${&�W�~������Bs��4"�+}x���`�^�fj�n�e�sc	1��TɑS�.�f��6GT\��\�,0��2�~�yV-2� �{�`R0^���w�"��?Yˉ�����k���,�Iá������\j��1gMJ����M��n�d�a1zS�@��.�i
�Qr�XX�^��GӴ�Ww��!��'�J�Z���H�i�?��^�풮��ݙf���F�)��c�$� �qZ]�=�u �t-)	΃$��a)��#ʧ��M����Ts�,�q8t	�<���ɗ��+>��|�^�����,�6�X�ì�N�Cq�[�p���G��{>��ND�(�����^�&��Ş�{4X��/�F�,?�$���<O.w��y��;L��2��qa���:ƚP|~�G�����i�����k�3y~�����*���>�Y�Tŉ�B���C�78<G>�#�75�4Eo9S��4	Ռs�_}3g3�E�����m����ݨ1

��}�M\�=�)	]+���-3����]�}��L+�BC�8¨��#������~(LF�|0Yq�(����/��7N[��L��V�z}�e3�OS�A�Q�c8n�	V����Lc��3�O�MRH7��A�S�Y"ȿb�H!0�1ƲX8OeM^O̚ʗ�x3g��J:\xb,]�1S8�c�`�Z�K�Ŝ��*�7� c�  9$J������-�\df���BD;/�-��/}N�R�}A�jN(��� �z��v�@{��l���DJfw�=B�V'��g�'��sI�%ya ؤ�3�Cۛ-i�x�x�o�-�����5mfN��8�<�S�N����wIg�=�7�=0ƂF�Í��C�Kta�<�jl�*���yf���v�q�+é��rǲ.�hۮI��9���Y��>�4p	 1om��"�G�����O�$�M6{���.�;�����:mu�c&�Rũ��g��e���)y�	�>[e���Q9�nS���I��B`o��r��~k@w��[,P����zע�"�1��;b��>���~r��ug�[��p�ˡF�6b�_�z�8�a���u���3W���S��*�	�/����+�x�������Y��<ء�#n�,��<����{���d�ݬ&��Qd0�U��`�#0�g�G��d�%����JC�:����Z��߰ImI�	��V��������!�z�ˮ6��Q(������Ye��6�ã��6�D���>�N)�1?FOǦ�Pqxyp��^I	�bE�$7��:Үi�؆�R������Gx��do�;���L9�r�&Lx�0
�#��eą2U�`���g��;�ތ�z�o)1�t4q�T7!Zl�1]|�GA��K���C�E��_r�e �������u�x$�\�7���py2��� ���pR`�K��x�����'���.a��0�bӰ�%��X���0WH�ZG6w��STb�F�S���~�@I���=�x���@��l��XD+�$>֋+�^����H����f��\)@-��0;�^������*�]���C@���e�฽���vh8��5�x�`��o`4n{�:eE�4�,G�"���؁�Zܫ��Wuw��ɸٙE#;Ո+P��<O7���b�
\UV�C�:c��T�7���:�{C��7_�:��D|����C��E��6&f���_����Zz��?���P
�v���1
t�Eh{�GZ%��]ҠA$�c�ر��],x�jP!��+}��ݨЙeM��T��9!�#my�5��m�O-�[ueU:<ekԺ�ke+�%veh��0�-{�j�{��]���ͪ���"Q{ާ���4x�F3���5yrI���-�K0P}"�j����
������`G�-:�K^��,
�۪��
��y20�G�����!?�
���q�(�.k��us#������s.����g}�f���]�H��:�y3��Ԕj̻��/�p�{�q:�!�L��K�U[4�Bgϭq�M�W�2ڴ?���9���fwJ�"AD�0��0Ć���iA��'��'��]���FΠ��]T�QQ�r�����4�`�Iو��Th0�4[F�ᣊ�.ǉ.N��O*QJ��?��o�C?v�+4w�#��U�k����՟t��Ӓs�j�uC����}��&��R��7�i�Պ>�s�n~H�A�����N�0�q�u�dw;>����&��;束A��@59WZo�y��ci �աԎE�){���-�(�ԟ��s�PEZ�p�$���냋��ܻ��M{����v�d
��D�8k��+۪'d��o�W��hҟ����#�2�1$x�� �FL8��k���}�sI��W� VA��#8�Bv�	�s�-��b��A����B[���о�ht ���#!%������-a��yc�P�8��Ǡ�q��O��Ze�,�VJ� ]���78lMc��m�ɜTQ���{�xƧ4G�3�>����}���j�������֙9�

=�J�Y��g]����8,���豭�v4���Y�{���������]f�N'�k��߷[D�D����d�o����%��ּ\�h��)��B;�Y4܋��T^���u{��@����wv(>�Nu-J �H��>5�m������w-�
|G���ɛS��n�3��ݍ�N�@ ~�|��Fx�*��:G=���.��Q@Wƾ���6˫�'�"(um �`�Y�كNڏ����gҊ\%��� ��S��?�`N.���ěD�^�.�T�a���8��,`�7�e��Z*�t��}:<:;��:)h֗�12�V�2����Y��5��\�a���ߏ�k%��w���z��������t��O�9�=HE����Rx�#�*�Aシ��o.�od����2�"?�F��(��Թ��s܊��0���d�U�H�w�V�_bq�7çڄh��s-����s8��Aұ���Y��g(��eL	��pۭ�=��`A��c���Y���ۡ�����]���;`^o�K��2�Y�ޑ(�(���=uxЄ��'�.�#�b���+Y�q���~���_�����#��f;L'�H��l�^����'+Øy�G�-�U�,o��c���-q�(��L<S�s!)�A0N��Za#��W��|��7�4^L��4�SXXF�ڦS��,�2��՘���9F���Y����빌�?E������I��Gd����c��U�7g��F�D�꽘�'�]Џ�,�gR���{c<A,wk��sG�^>�կ$RA\�q2� �+_ǽ�V6����!P�R��2$�+�wX���$6�m�I���٨<sL��;��=7�I��L��:}�gj�z��X�䣦	�pW͵9� &�sǈ'��xq����[(#\^��{8Үr
��"�;��"F���oJ���Q��,+"V����v�J��ͷs�'!�~��i=�A��6=d���[�>��y�,i��2�H�F�XA��~Ttc�'���Y_�VQ�<Q��>��A@?m�/��
U����!�{�t�U��[���!����S��_�Q���LM� $�7	�4p�HB�!W�ì���������=$��S>-W�.	��$5�m�r��2�S{i�Փ�U����1j��v��n�%?�]ѩP5l �N���vc��_h�H�b��etj����{1�)1&�M�	�6�6�C1���~�����$�[1�m���uq�n��n����;Xq���@�Eڻ���P��$M@����b�@���l�B�769�JCa7���������n��$id��d`���Z���b#���~ΆE���o9_L󀓞����`���/ksZ���|��	i�-��8k(�\ U���;V����7GMLh�Y���|��=o zK�O�jU�k� #=�;1J��o�c[��*8��+��wM\����P�P#@�2���v;;Y�G4I�YVMB�nr�� qg-rr��'m=l����Nu~�(����Rg�JS�wP�Vy��"�o��8�������m\�mXgV�CL��v����^m
0����T��9qN��BE���&�u����~��u�'ǎ��Q¿a]��!�"��i�X� ��~_�{-�h�����-��'ʈSC���tc�Շ�r���r�b3 l+��P�;�4p��-w�^�=�Zk�2h���i�i�Ůi�1,&�����p?�
U�����a��i(�j�`�����A��`p1�ik�Ū�Cx�^"�E�VZyFSJȣ�v[�)	��0�P��8� �`.�L|3��;�B�X�����F��Qi�XRߩO�Y�BͪH��㮉�^� $N]nM��um���C&N�)"r9/6���|>�����N�6W�X�Q�_��Hd���it�y���tey��ѵ�^Y�v��l��A���Y=pΒ�v���#My8�*�tQ��>&����x8�-u$p%N��^GL�V:[�NB�~�����Gx��&^h7�YDU��=�8ک��E"O6ʨw�,�ϓ�S�8����wO�_%a��L���F�Z}�ҤƄ(�p�A.�����)�y|H?��^���_.�'tU1
�v�H=�az����}�n���\��R0���&�Z���L�NTߑ<V`��p��5yg��vN�k��U�Y�jڅw}3�Da��e	�+M��%G������M.>�D�dc��D��c;O�Ëd�jD�/�"��δz򦆧R�� p(�������m�簱mf����đl	�eO0��΢��W��]p}���/�6;A���@L���>�iԾ��L^C��@$o:�o�V��]-g,Лz��v��ad��!�_,tw�J��e��m�����Il�E��e�n"��{TOr#�Ԣ8��S )�`����-���Q�>�So����Z�H�p�D�q��t�$#v.�	ph�_�F�Y�*����%�E9�٘�:c�遦����.uz�y��@-�霑�& ,y&�PD��Ά��2�w�)��m5��2a{^c��Dȏ8�P�@{�d G�:'��a=��nR�<��erж����x�|TAM>����B:ć�u�ȓI��J`�Ka�-$@c��+��m����gb��H����듒H��0���lnΚ�Q�DͶ�����}"C���jI�Ld��W�q����ն����MzE90��1�N^�~�\o3�QK���x�/	���k�u+5�L"en	~Q��d/�J[bˇ����iaoEz+�����-�	��]�����i��	d��[�Z��m;꜌�ɢzGHX�(�@.�}�`$�~f�/,E7��ë��dj��'EO��}����
k��� F&�?^Hp�&��Jg��'tV��:���(�f��5�3*%�hZ��D��
�=��ð#� �CL��ҌC�pK,�M.�q-؎��̼"�.^�,Q�0�m�Z:�khk�x�;f�J��^Y{�y�V68������^��rY�(�d�g��
�R!����|�Ԡ]��Z�H�k����O��w�+��6j�	���@�9��/�K��}���"��(��3MgЏ�v=��f� ����ʡ�{�b��a4�1������H̒�iԦ��d+w�0���v�����JF�G�0�����)f��!�<T%��ƭ+�bPP2(��C�+����5'	�O�yc�t���hz�r��9�r�o����[�&2��='�'\p�Ԭ�z���1n����<� �<Z����h�]k��`p���i�g�ݶ�7V�����J'2�Y0en�ȧ�!��޹F�5�Stf[��z�_��ܥ���1j���=�$s_1�ZKf�6H�=X�8:=�U&q����ώ�{_�A�o9Y煼g]+�*�Ή�$��;�؄�p*-�U�DG�������W�[�;#7䆘epg���)j�ؐ#f��I:�^+�$E3US�fYפ,�+B2��[��"=a���BD@�`ohf�0#��5�\y~鿉�E��in:����ո����wҺ��;-@P��]��-��dhu޳1f+��]伏�Y�ĩ��xJ�ʙ6ތ����E����������g���(㸨gu�$ߚ�/�t�����uY7�Pk�5��ΰ\��'$����*(ރ�!�N6(vL�!g��w_�$?l���b���}ϡ'<:^����o�xK}��L�$�엎	]2��s�����X˪To�vs�(A���)�[�q�yRjy�q��/�Á�*�:�`�<���\�3�A�����U���C��0��e�`�
[��`��U�`N*�5�7�\�ܟϙ�Y��]�$���������g���^�$��;���7���ب��R��[#[��$K	��:ezf��S�]@5aC��
�K���a4*�D,��ʎG��_n�B�3uY�;^�#j`���@~e������FXi���ꔵ/c{��B����4�y��Y¿�-n5��i�"�/9~���p��A==��P]���nMC��)Z+AR������0��d<����s�>��a�iLE.�����4�'���.�E���b��|��:�M3��f�T`.
���q]co��fɎOQ�aӹg�)��<|�-	�	Ƅ,Q�d"9����>�1�G���~���`j��}#9Sp���`�}���n����#60����������(g��h�.@\ӏV��5������v��P8y�o�������Y �<��u#B$Zq�	���cز`�����q���9)?٭,�&��+iziq��7c�x���5��w��e�8�=�`#l��/�)�@�#� ���'�rJ(�+�6�dg�d�O}�t�p�Z��`T�ZP3� f ��ӓ�T��qm��^�@3�M�2�Pލ�
eQ6N��Y'������H�H-2�t�(��M��h�]&�ٵ�2��r�yA$�{G��>���ă��k�'Ĳsc&t���:��s#|fɮR��1�j(T�^���u��P��ax��r�#L� [�%�-R����Hb�l��"P%�Ø�6�c�i"4������!�$��������*|2|f�}���_Jۼ'{��`_[>�9#ؓ��k$�XG��H�<�L�LH���{��p|)�6]�';�.�"��^ah��	:�^��	)k�g�{!:B���S�$�/Z�&�r|�����.��67�I7�Y͓ة�\s�Y�jٖ�'B�]6xY��r��]�Xd$T�s-hb�Nk��$���JP�9
֤�c\g�;�q�>k��e����~pn�KBbgx�>��&�2��_��-c@\h�_���[���هr]Cx�%\�[x�l�t�}̮f��孨Tk��:�1���ϊp�1�q#��9����G�3�D~+�<�؆�?kR���r{�P�7#���ɡ�|����+������Hڑ����0������w�p� J3b"&z�ͧ�m�|�|3D��,F/E�_��d�se,�a�+�`A;&�[��TD"��OcN�eb�K�Ld�ݠ��_�O��n���z�U�/���0�v�Jc��[;t3�AT�u�ܽv��8Q�w+��R�fCD�4����Ք�h��%��`�e��o:6��(���A�"��S���sl�(ZߧB-�\���#6sv��5GQ �Y��*F�ܑ�
�OO�X�� �<���5�r�5Ɠ�R�5�lW<�ē"#JR��^,?�Qh��\<o&xt�����?�-q�$7�+�A����a��]�w��J_-m����?���|%F��Y�0�KX��n�_��A�����ё��Uwc�cx��!����Sy������W8]��R�A�+��ɹp6���t����s��<�%�#���Жg"��U���#△�������p�O��6�~0c����-��6�ǺS�%/����n�$7�=�b+��D>��M�m���Pǘ�+=s,�x7:�8�(�b�4�r��'�X���i�-f� ���zZ�
�]�A� �R����ܱFo�|��&�BHO����^��fCs=`�{h@�I��)�����l�Ƕz*����hS�H��LϺ/����1�琫���faA���ȕ��t?e��#�#�e,�UgD�+O2lf�0�����Yy#,�_�R�����4lK��~)$$�G��7��&��1����eFL1�Z}�����^�=@�T� Q{�栩��9�qh�+q�6'4��ɵ�Y\Μ6�4��Of;�KzF�D����#�b�~��{PI:%
T�̤�ʛ�Hb��q��e���y=�����Ly�/C��L+�����������{�.��Xv�ӄ�į�).H�P�7hA��	n�?0~��(�+�����m�jf�7I?�kxZW#�D�q�%�������=�����K�N��v;��}+�=�8Z���'jv�9؃��q4z�A]�F��x��&3��-�o��yJa\[:��9.��z�����Ӈ�����`K}�.�lG��=�$� )��ˡ�FV0��鬬(Zp>�״���Ԩ���_7���*��7"��xohp�SǕ��j�jϚ�i�w5�oN�J��&��?��
���O5a_�6R#�����7�T5���h������p�Rѡ+���j�v�2
����.G�5�u���{�Ho��~P�z����S᷄�/YF�:�ji�}�{�0xiP������=�Ԏ�WZ�g_�Zݸ�".ѥ�Q����	z�>�}�cO�ҭ��w#2F>�
pYي�:+�	��cb���^���x���	�:�|���\�!�^�7��H�F"Zgh���0��������7�}T��EZ�n׏��:?�GQ�Z�ǚgU '"ߚ��=�:��CS��Gbg���8j�	$*뉞�z<b���I���`b�S�̑HT��n�$�B��G��'S;��!l>��$��R^�)��s����.~s�^k1H���N���p֋v��P3S�ՙO.*���7�<
�z���F�Fە�L�+��s��g�@P?}�J�o��<,AS`;�$�Ŕ݌9��!�p�5o��R��D~�31m���B
����a2����M���X`�S����d�q��Fڑ7�`�1�1�6q�'�$Y֠xZV%*膳��� ̲UPeu�-�GR�>4��a5
Yo8�=[m�4�Q�����|�!k�k�Dր�繈S�S݆e�������\�4��(Q�6�^���� ���,�[�<&�}+�m��64X��a'}�_|����(Pe�1���Оn	�p(��:e�"u�a�ϕ�ЉyB5�N������g�i _��y#��p��募Щ�d{8��2׏/�70Xݹ�_J�*��V`k��y~�[eb��n�;#K����-��D©�p���|�ϦR�=]�_�l=q��ô��-}ĩ`����$Z�b#jNi�Q+?��W3žIA�)����B$!ؙczf������A�
7w��Pӷ$�bƉ�����A4��-_�$~�h'g2�.:�b��o���U%5$6ݤ�f���k�س(풒�fR?vY����L�}qB���mAG~S��]@�l#6�㾠�={�`�Hͪޛ�[�����q�Y]�XI�A�G?޸�*Q�m�:���8�g�D��X%6I�J�,0� �Rڝ� 5��b-�69f[�5��&�2�_�,��H|��L) {�od�D>
�7Cj'�������/ڀ�t_�1S�+q��n����c�E�vx&�)�x�+�X^@�.�l]������7���W7~v��VP�q�I�
�Z�n��c~�Fys��� �&BSf�	&��U���H����]��>���rB+���mqJ�f��޸��3J��7�Դ-���|-�J}��T�H�N��gW;�$��10���64�����t
���p�&G���K@���'U��KZ����Y4�^�Ku@�Ab|�V+&���i���#(5�}h����IG�S��|LC>�<�6W�^$�9B���4������ zn���6$Hf��lg_�<ܺ�r�1�en�<�=�C�ж� rg�'��gW���ƈ�07�]���T�$������4��ؠ�&���i7�J��g����F9��4����r������=��Nr%��49�<P�@VS���e����?Yɣ�~\O�&}3M3� ��hsl�1� ����O,��-���z���P���=Ж���W��i�{���q�gԏA|	>H����U�8Hgix\�0@����'���ko��7hӽ��.kD��mgF0���*�lE���A �o��p�m�dC[�@�s�&��
�ud���K}� ��_�0r�xD<h�rt,�WF'�e�NY�f��M� �ڂ�/�@Y���w~�\���qw�xE���`����H�@7<��A85syK��,Gz&�� ��ZW��~�`!�Ge��D�[���D&z���1 %�kfY��<t�B`JR�u�¼�V
��o�w�J"K���=2:���:f�%$�:U��\���d�"����?�&��@�����HY�F�S��B��hS�]IKS��M��/�;ߦ7_�^�LԌ*V� �bp�Ӽp^���n�
dC�g3��~���Kg�p�j��Xc��o%\�2�3S�*���	-�Ϝ^f����w3�4z�Z��7�*V�gR� C����g��J��������P%�[`hoY��ˆǲu$�����/��a�yxOmn�.�Ƽߔ�ZHk-XBp��{^�Q {	݅�U*���w:���7N7���_>����rh!�{S��E��� '��i�����L8�́#5����gfV:i��2Fq�{���׬��^��o�N�Ȭ��v�Up������\����*�,qW�3�ب�q�z��23��w�����a���3f%֊5+j�,{^[���K9m�3R�^b0Q�o�5H%��Q�
�܋�_��y������U���}�Pz^;�V-v1M���,����G��D蟔)�Z�z\j�B���$m΍%�ݜϪ]@x�m4J�u�ѳ?���P�7!�?e�� ��LM�vgh�B���U���Š �u8m� cGb�N�Y�ߔ�!B�3;��g����;�8[ شƗh�2�@�yt3�~�,i#�}y���*m�i(�v����>LԃD#���Z^69�O�]+4)��Z�F�̬�`i���S�����;�0;RcB*�{�یm��Po$��+��8dk��vfQ�T�j?mr}ߪ8�e;�>�ܪ�Z���i��<v�r����pO%�4Y�Tj��
"X��4���,:aL�������Hᓙ�+�c���fgᘤ?�?��t�qi$e������\i�_�wy��\�w��M �SEcQ�Q��M�{cBx��&�Ƶ�F��\�4�@�,��&��F�o>��a����}s��N]�G0�S�� �Yoֱ��
��R��|8i6�xoaO�>H`�ߓ�q!�B�kH��>n#4nE(4xk|���CR�'���"����UL87/��*���bf�Ղ'?�R�&����%�����2a��c[�$�e��h�!���۽C+w��y�3�O�c�����сk:�N�������I���ɪ:d�4�o���G/=W4��;*呁�����vr��OF&�i-�����Ի$X���=�_c-�-K�]�A��G��ӗ���7��Œ?�i�w5�`WK}�-$�t���[X$�� 1Ba��.����ּT����M�p���Sބ ��D�clho������^|��#��r��YC�f���C��Oa�v�dk����A�����l	���ڨ)��`O(=��� �6�z���s�]���|`K啞>gNtq�xa�~����t�����Zb :#�}j���yN�ؼ4�����6�ݨ���B��$�Ӳԧs�Q%�2%$z�����ʋ���rƧ��<2�Wy+�@`G����!�,t��lX�.Pkæ��=]aO^2�����U/�_ir�1�r���7�gY�����Dl��*��(����r:Xޡf-(Q��]'�ȓ(FO�4b\�:�*���.�|������k�I-�^i����{B���*�;ĢJ�6�W}���YN�,�1���{V!ZQ_�XR�X�JZ��ZR��Z����c�`)�+5�:���(����O�=T`�i����e�������@��b�R)	K�?	�-���(n���
#,�0:�"��CL�N�-�W��!���C� �P����s��I��H�?��/�U+�l�OQσ��������(��o�.z�T���0b�!b��s��m�x�����L���DR� ��Ya��U��kj�D��MɆ)<0+�D��m֨����Oc69%t|�/mu:�[���$���T�gS��9![�����[���0<u�����Zj5_c�d��+絟����Q�i��!��0��3V|�+���~[E�M ;=�Q+t�R�Z4P|
�2��hƘt����u�_]��!H7!,�x�y��J񚓧��1D;Z����#�4fq��"�Ő������XC� 0R��<��8."_�|9g���
����c_�c̳�&�ZϤ���+Oۙ�ӛ��!T'��nI��g��W�����x�*����mR�*z�'X�Y�բY����N�k�ц����^�0�`��*	h�{ݽ��T?������~�ͬş��U�;&a'f7�ݦ_i���K�������$���R�~^M�Q����@e%b����z��`KV��$ONmw�.fVm���$9+�V|L��c�q�N�e�����Rx��G������\��(p}�z&f 	Gw��hm�G_��ZR�|*#�ro~��͛���|)&���.1G�L�(6ز�^�R��u8�<���=,>T�7)�5~8�wu�6��i�դ�����$��y������kEH���N�����������5J�P�����j�:���H �SH���[}.�fq۶wI���cg�wl�9o%V�J�~�
�����è����,��+�v�`���:� �;���s1$��u�����Q'�]&�em^��aU���z�"��!���JJ��b��D�ȼR���#��4�N'�y:��^U#�"j���#�"Թ���L~���r��	C�2�KG�,p�箂��ܢ���x"+��������Q�-��"'V��?�#φ��ħ�v$������R[����c}�X$��^n]J��ҳ�J�J�P��?����S9o<X� @�2pX�u�����I��Rv�p�9F�O����J��F�C��{��nUG�Ku��JKA.ʌy�7?Q���y9�8TD7�7Y��"1d��;�^�����e�������,~X��t��9��D2�,GJ��9�����!�u�<ly�'��`�F�P�R�f�\.g��GU*vq��U�D����\4X��au��[�����]�Y�o\v��]�k�(�i|��!��c����	��sܬ&!��8�J9-G�-�c� AN}�w &w�Wg7`iAH������J��P��5N��y=��8
ǌIB|%!����аx�Wι�"3R}�����sk��,j���tf�_����_P�!8���d�y1����:Me���!H{.�A��E]��ƍn�n���V�����%GK��u�P3⊩���Ý$�������~&�h飪2�01���	�>�'<qz�==)�͢�]�?��O��|B� ���n&�͗���\.���ߋ�]wM,���n�(���&�]�������U�T��[���������{�B��>$)6i���ih���7��SUfV�](u>�E�m@��d�p�i�>Z%��%� �P�v�(��\��Mg�L����L)��TER��t1P�̾Pwo$%)� �� ��"ٌ��m
vOߦ���Ηf��p��F/5s֞�$�ۺ����P7�����̿�]g�18�+��,�b屎Pl7:(�o�-�$ߥ��O��+����`�T�_'�����&)��"�7��G�]�����R��8�Sn�2Y3�"����_�'/(iͫ�e�o��tZ�p��X��\�g"G�V���M�Ў�2�3�%C��?�ϰ(^y����4I3ZH��6A�fU�Q�t$����F6h�5�i1y�} 9컳0��;*�
'������w"������*WZ��W�wQ��͗�����D��F��d_Cn��q�qi+��a������Cn�Չ�M��n�MN�N_nY��8#I��/	�\S#\�N���R=��HA��a�G�)L��E�����}+~�w
O�q���l���B�s�P�*����`�)��@ƨOĉ�l�imߙ9j�5�!9���4H#���mm�M��#����$�����x�@
��Q�FZ6��H���oG"��O` ��C�,{�G��^���38\�ϗ�]��pA��}�	��^$v��b���B��k$,���V?�4D�]�����sLv�h���o$���t�~��ÐM�b�.[��3V-��OM�{��<H��?���C��)���W��?��F�z��j�z5�K ���>ؐ�5�	Ez^�t�z�׹�	V)�aZV��@G$W�,��^)�*���/e��4���<V-��/~wt3��A��b&�
Qa�0&�K{��/׼�EM�Z�G��]u��S�������E�"?,�أ	Up�*�n0�-�1y����T�G:���x�Oz)=����_!\C'�I�����5C�j��e���>�����mC��ǽ��z�)�I]I�
n�!$HӺYT�՘O�,�a�O2!�Wȃ<Y�G����u�,RY�zUA�㶃i���Z�{0"$uC��▪&@�qM5��yDU�,������=�G�gp�b�`x6E�U:>I��t����6����/	�OU������k��y��@ËEid�fO�BzT��湖�^���!�~R���Ô��9���d��n�(ݯհdQ#����!����θ@��!x���(} )�ԃ, 8��%��6���+��a��� ,��ۂ\�{�y��R0n��bm�F�_)�,KWٶG�d�1l�9�Cޜn\�R�D��Рֻ�(}�9$w?B�����M ò���Y�*h �]�W^ˑf�w���	��}Z�P
9+P%z���v��X7|\��I���'�yT]՟��hD����< �}J�T	9�9͔~+��YѯH��@8��r��Կ�(Q!��A�1�����R�z�"�S����o�(v���R�������?s�d�'��Y�yz{*1xy��(K"�q|��Vm��8���D�jӥ�K�_~ɑ{�<�M��}���?��#}�1�6/���@"��Q�$��֊��b��2�,ԤP��p{� �s��}��K�^������;���į�	�n8��^~����7�a����&���GKl�����w��S��7�ί0���F��|=���s��QɅ[�����f�J�������k*�3֌��O,m��ߡ��?�b?�6��v��P�
!�1�o���g�f����Y��Ͳp���8(�
��KC�����M2f7ɛ��2�b��@���u�p�� ����d���Or��JL�bm�����֬{�c�T�\�Ђ�Eo��'�B��Q_��s6��顄s�v]�<����t{���AJ���u�����oSʔ<�o�a�?<��~�5>�6l'�3�]�an2cv��dc��e�{c��-xF���
C�q�J�m��/v
|���/}��*_��zÌi��1�3��K�kM̉­��zR ���2�q_�mp
�ba���Y
>�Y���$ᤄ�|j��s��_@>]KZ8*�����n�i{}��1��B�Ob�����K�8&��֋2��;Z�bG	��Ζ�w�]��N.�]@�w1?T�������VX�;�8��� `��{sY��HV�+�p��jga�g�T*�������*~EO����\�����n,%h���/ǿx�X��������]=����W�Ua��Q�7�Z�J�p���"�����$Q�4:�<��p�r;���5T�����	s��ٵ�#��.�j����lR�D4I��3T��~J�:�c���/���!�_��)�!�6����1�g�`�+ci$�߱�i[t���x���_*ܥ
��n�q��^��y�jVO5��D�x���w�89��ugQb�x
�%�(Y?
���܉`���:Yi����s�y�?ů֛���l�N@.X$GѮ\&�JZټ�6���;v������� �Hg��9�f�w���\���)�u�2���i�+L��Y3����Ž!���ZMT�z2���|�3|�/�u����P�<�J�9�oi2ڈW>z��CoYz��/�l-� ��\���!�K�H&�8Jj�>��!0�:�씰Õ�$���> �l��8^ʄ~���ق��Or�>$%ԍY�'��?��L6V�j���D��9~��w���J��G�(��s�p�i�
��B�ބ��i]}^�yj��rs����x%���]�5�$J��b��7
q\��KN[Q�S�"�ᔳ�m)<����JK.\FA(�����)������<�(#w��?gQm@�b�*}vƭ�>/!�y���^�M�^����r�Fxt�4ﶉ��)��ӷ2%Ul��ˉ���)(���Lغ�/f�au��Hu;�OTI�:pO�A�U�X�ǆ����b��s���Y��r�xNO����j��$�����ۢ��~z��Ҥ��g��a Cݖ)�# ��F���,����/���MA�\,z̠�/�v<&=BjM�-lh��M����B&XG�@]�	�`���,d 3�	%⼞0қ������W���J/#�vM�Z\a�&d$��>���c��+��q�xM�
hk�,0����z�?�!�9hm�W��;&MX(1d��L�թ�� �C`�w	�/��|&#n����LxPt���o�V:|��b�h9t�3S$EE�i.CN m�; 떈��$F-e���8�砵a!gŁ=#��׳ aR��Y-4�d;�S\�8ZV��܁Dg7w&@SJZ�����dU}�-<��!��LO��A�M�#��|��jq��k�^w���/C2���x�u�Pj �N�����^�NeW��щ�Y`��o#��ag6)����q�M.G0����%��/��v(��ez�.��?�j�W��ݧ��<���Vv���1��bl*�kǣu\5����g��d� \�,-G�����QƆϯ��ڷYx��b9;���:���ch��0�Ta�;�Ң0����ء����z"3�*S��)�鄶�oU_`nL�{/N�]ߋ���˿�I4s�G�eڗ8k�p� Nf|+MY�I�ԴI�G8��Z��I�BIw���|&�Ĳ'��Ū�d[/KP�^������� R��$8�Ѓ�2l�7aS��J�X��(&�U����/L�p�t��&�f��LS&sEe�稁ֵx�1��M���ۖ�WZ�	0�����1z����?K��O�S$dg#�Y�lxj���B���R��G#�&s=i_#Яy���.�0(��Q�#��g�\����w�:з�[�V�@A���	Y�?4]IY�����Xu-�����wV��|�}#��g���-��g�g�L+m�`s�"�k+{��;WB&s���nN�����K�gJk��^�LI���+ 5�<�D���!w�b�x�y�t\����{L��*.��X��9��ki�e��_k����S�!�H�*��jLk~%��'M����3pH��� �X7��	����ko��@���?�i2'���ŝX�XdZ|��R|H�����>[��~���t���ċ;�Bݨ�����J�G®A0[��o#B�INi��_�,���L1]E���=�$}�N��?B�yZt�VB�y)���K�d�������w6�)�M��MY��	s��%��&@��rb�^���E���ܫ�b���Y%O=���h�����"(k0>���6���n8d�]˙F��*��SB��7�%H��M,)Y��R^v�f
�π�H&W�*W�P�͌�q����R���F8\E�1����.&͛^�����]>�Z��9�h2�Z�:�wΗM��΅ji�}�5�~��[�����q�N\�
�4L�����ʩJV gk�R�љd_S����Պ�z���FƆ�8B39pF0�S�2rr��ۃG>����>�x-d��n�nZ��dl�>}#S@�n];�[�ɴ��8m��!�LD���4�yE��D��f�o�ŚVR�D?l��ip:���b-���)�}����)�$�l��p�1&��/�!T��)�<|ت$ɶ�j������p�����y7�p���m���5Ė�H�3�*���H���xD��"N�1AFW�)�[�_�e4��&����dx�)����҆XX_׀S6� �
�d��<���jn�M�{�v����������$�oC^g�y8z>�&c���=��_ț��z�P���B�ȓ���g|䅋�_��7�%i+�fJ��K��RW���YV`]�&O��Dŝ��&t7á�>�u�$C?c����0�t�I��R�d��͢��-
���LU�E��w��
��!��Ù���c]�>Ff�t=a}\�G�42N��z|�ix�������c"��K��Ѳ[h�A����"�q*[

u]�%\�X��Q��|�Z;��x$�;�^(n��u`f���Ɔ���"���ɯ	�w�a�QMVӢ�5#�@`A����A�ʲ�,ZX�N����(ط�^�k�r2�9��o^�|f&��kZ1�SJ�ݧ`̻��ɂ+XQ�X���DA����5%�ΊK��!.�ϩ�vV���&$9|�?W�=�y	K�|�W��YR
�v�`͂�LrTaJ0�/�ߚ4|�O`,�B*���Q&�(\�'�v�uSdge���(�V.�Sn��2��**)�&��,qx.�&L���֘3+y��#MS�ײ��\E�2�@e�7��DD{3G�=��IB�|D)��+�hi��c�c?�˿�J�!�2�ٳ�A��j�MJ�Q�\�G�s��Ŏ��u���1�?t�P����W�o�?��ۿ���?��4�YU��''n�y�$����!b��<J5jo�~�H��������ީ�vi�-������Ã�~$���'O9ݜCp�y�U;�@&�����*�dm:@�zj�W�Ux���,Ev�EZBj��zI45Bq�4����7�+�%��4�	�X0�D@7�1��_��[��]dv._~����7�}&
w)i�B�3d8G�\K�w���R�i����H3\7./�2?�;j��}Q�"~d�(Q��������GȀt+��24�dЭMs�w�Gڍs�g���k�-d|��^B�}�Q$��p�U�&ڼ����[�]�t�?$�%��@��%3��^̡(����؃��ۑ���o]�&�v�蠗�=+
%��<96Jj��i��#����F�����N���}��WJyȥ[���~
e�&ՙ:T��]�k�#^�af;��$M��lh�ff�M�X4���Ywy�8��N��0���S���;�I�G���~E����f��3l��4����J�`5SsY���-�YzS��(�
�1������H�͋j�IY��d{��<`܈è�����Y}���?'�.[����"Q$e�!ZX�����wD2n(����*��gUJq��;�&�3�X��t����ok��/�G�N���dw�t~4�����P6h���������$A#>�F��RH���M̻`�]c��o�f)��[��X�me��a�<%���J�~fX���Cqǣ�'�>w�v�$���cpC0�kE=9Ocf��]����2�����Dy	}{3�[ә�R.�;��w3,"��L�6U�ڢ�q�k:D��lQ��4�J��%2T<^�Lg��M������y�hjx(;�YR� \��+�����L��������Q�s�"Pl�k�2ñ_���.��j�G����xZ�ψ�Y��!�O���Ւ$^������v{�	X`6�mN*}�`W�\f�lRQq�(`�e�2���U�ʵ��)yO~t�d/��ٞɌsw���VE���o��%P�25PE�S�W��I�lY�����A�	����$�E�R
 A��o�~{*�OqX�e��++�S�xԱ��rb_Xj1u4� |����p�3�MDv��Ym�a�����<2����\^T��ƮO&r�/��{�\����pG�h�z���O�=�|ƤU����Z��2"��u���,'�X���5樉��W�vα�M��{�£r�x�:���P����ye�Q�B��͖M*�o8.�;=�u�U�.�h��q]��&�?&�*,��,���V̇eOh?Ϟ���gT�@�4��
p9D>U�c?��{{��4j ����"��R��ztP��Ƥ���>
K]�l�E+g�\E��G;���(����킜,��'YW�����D=H�&R��.H_���Ǝ�-���۰��+�w��wm�gcp3������ѠN�&|*��N�X,j:����@� ��O(Ա �G��V���!�蝫j��'�r�ى�xw	�35(���=,�G=�Þ���t��]N/����ԷW��d#��g����s$|�D�9kHRL���υFd��U#���P����)!��׽S�1�sn(�u0���a�Z�Ů��Yb�P���������F���`�E�rWo��?n�xTѲ�?�>��ARn������0��	T��
5g#ʎk�1�(L�<L�S���v�ĨD3�r�ٹ��o�R��M<�hY��}�Wx�`�K(���>��s˘��m������g�V��l�c~&��q�s����F�-Wʹ�/�8Q��
��E�G����D�i�p����h![܈K���,�2���=:�4l'cL=5Ҝ�?�Hc�d~1R��Uo{���Bܯ8�d���ZB�fMF��c�kL��@��^�Bc�]��{)�$=zց��9fL�-��x�Ox�5���l�,)g����1�c��6~H]��S����ɁK&�c��X���XLC�P�P���Sq"�j�!�~��$�|}�I�����e�\��9��&��jo�ٵ�
������5��FT ��dfm��1%�$�s0���ҿ-JQgh�kz�pBm�^��F���(=Am����6^l*	A���r:ۑ`=?�?��0�G2`N�m �8�4%���s�j�@�T�f��,L�y3�	r�rK�2�{�G�̘���}a瀬����=�Z��TԤ*+b���>v��߯n���w��v��\#��۳G���ϊ�ur�QWn���-u��r
+�ힺ�xW���zi� ���\5�s򰪤�J�tw��+:^��3��mQ� ���^��EͥJT��a�-�7��l�A|��M�>�t�>�&U}�I�),��x�iF����ѳ�߰�d���+4"G�41.1NO1��2j[�ɐ>�ϋ�1M��=K.`��lZ�`�y[��9��MN��S��"�a�F�o�ހd�j�"�/F-jbI�RK��ݬ	-|t��M
O��X=��SI�񁶃;4��x��]�,A���͘���@S�� C�)Y���wƆho�Ǩa�'e�F`%\�]��2/�������4�x���E.��	�n����Y��k��ng�Xa�H�<�ւz�ۜۯ�,��<�ϘcwO�M� g��1�:ʍ�Z^)�ʹ��y��m&3�zB������^ևF�,Ɔ"��L���#$r�8fY�
�&p칹�@����F�D	�8`��]t�k0U>)�Zh�VYE�ހ}���X���f^��?�6��w�����*z�x��Xb�l��\�J=� �mt�Tq�$|���7*<B�~�b�c���/��k_KP�c�����Y�՝}��) �)�W�~bF|)N�����I����2�w&=���5��wG�����7��pH�Q�85���b�U4-V* B����oa<��e��ܨ�|׳b�ٍ���Ni�8�����l e���䔕�~��]k,�*�(�>eto�ޝg΍a;�M�!Mmv�z�?�3!��j�l���ס���(ӽPr�b$��']�^b�Nt�;>��=�Js�fNS�9�|�LZ�A�w@Z~�� P��erb���d%#�D'���$Q&��G��Y�b��ũ��3*M�!�7�O���Kǳ��+�]M>�S�����L.g�	�p���&ϥES�*�g8�Fm�D����3�ہir�r��]7t.B,�;����cs�lM����D����^���e���p����JW�}.ۨ?j�G��\L��^�6��YX�ʼ�+}`5������Kk�q�U	��Աs%��s��
a�����Y5BO~R��&3�s��^�XʾQ7z�B�݄~� �oVLw���
N�$��>_ӄgs��Ά�0X��Jŵ�h�3��-��0������x-�̸�bl�7��m�T��v�H�PK���&D]�H*h��>zψ�!���
m��8�ȽD=
��B7k�N�}�h�E����+_a`�p�`��J�����P�DcL4��2��pV�\_٢�с�ܪ}H�7 �Ǔ{��mlX��������� 	Q�pi�F�g�v)3�� %ݧdmA}N$���y,�^Jr��l���~j�n��q�m�^���)�y{��Ѽ1k���c��vj�P�0�����4p�9ܿ�8oy�3�a���-����2�;hڸ��ϸի�s%okh��~Bico��v��:v�c�]o�](���$��{��a�Q�>�D�bsPn3�g���[A�	��u}��h��"!����y�Z0 �R�S�fփ��a3�Z�륑��3�IYO�����U��ݡ�_��ܖ�1k�a=��H&\d�(�~���"��vBa�����Ș��/dV��=���⎝7=׃z0�n���4��H�M�[ֽ{z�ͮ�8��|��U�k����Ŗl"OU �H�K}{��r'��M���fQk��ki�M�	(������6p����38p�&'�lIJ\���G�*� �8 �Qq��s??)$�e�xStk�<�l��®~��+3:F����>��?+��S�������"O��/�ӎ�u|��?�O�>z�oBS*�X��[�ſe8N`{��~�$�
�����%ڭ�CW���.�e�g������Iq/#u��������\�|DL
���舙������A�(�@�Ǵ��4��_�R�� �7�^�d��q�d!���I��e��5�+b"Qs#I�jG�H������?�N���):�*���q0�F��Z/;^VQY�L��P��3����F��7�[f�R?��A�R؅�������>l1W8XKq���،��UJ~:`!,�.�"�t�­�=�ߙcq��k~���5@����f�u�v��9:��W�����9dA�[�L��%4LH�����u^�WKh�ڌߎ�WK�'��),e>��=Vu����ZUZ�N�����Շ`���^<�ڽ|O��)�1�6岢De�ejlm��p�YmS0�'p8��vQa���'���>����!V�}W�P�vd����~L�+�qJ�&���`�y7��P����Ӕ\+4����3�r�z�>IS�u���p�ԥ�)�s�_������8t� ��p�P�$�~��GqYZ~�GP��2���~�W�� Xl�V<�V�t�^��8��C���F[u��n!���`�ϱ��Z�D�s_���R��}��(k��:���4{EK�n���c����f\��]���A��/��12w_m9K�(�����P�	1��x���J�q�����j�[2�JL��n]��Ա���Sq�!����ڞ��`����;����ͯaC��j�f^�:\�а	�]l���`�I^���})�>]�{��0$h$����#S�-��(od��=j�'��e���G�c +���un����}c1��7��tp�r9�_�I�����P	�pl $;c�g
$X���N�/�j�B��gѡ&�I$�Iu��P�y� )�ne,�����m���#��Ó��?�s�J��y;ut�nc���R26�l��)�	m}֝%�0zF[hD~��갷�~�4^1+ӹTC2)n?�C�'s���s{� � 	�g��f�܄LE�	��xS���3n�?�f�ƒ��Mң��Vr�|+��kX	3ԡ�ȆDX��#�gSV����z6��'cȻ*�% BUJ�'���t�*���RXY8��k^R�q�m�\tW�p ��KC�B��t��&=�@�ñ�:�[�V�L���������y�I!:h����vRaB`����f\I%�g�d�d2��Y��W�����2��̒cBe�'�vX*i�/�0�W����^�/�������R��2�=Y	��U��6u(G�)����mg�c3�w�UHWs���1ZJ��̈Ob��L�F���=a��"�R��BX�?��0O�6ޟ�jmF���f�X�K6W����l�6���.3���8�OL�c�ɑ![~�P�ep7Fze��"(6�l�:�e6�t:N@�Y4"&���j(��+�DkS��q�k�,�²���!���&�����y)[��g�
�e���̬0+=g���A��h�0���y�_w1cg<���S�;���4���ֿ;Y�-
&p
b���H���zTqR�|�Su<�B@L:^z��E���d��.�a����o��	\��0�R˰�4A���Y=7�;A����\ic�b�ۧ�n��b�3{?�ơ�VMK?�4=�0$�<_�ԟ?\q�Xǖ8���u��� �e���BLk_r�����|p�B����'.n��Z�� o�0�!�&D^4�38�'�HL����/1����E"��gg�<�r�����t���`7�/��7���.'��>�`=,���#�ώb��U"}�B`�ƛk����MR���A��6^���7�1�y�Q��o;7�����#�׸Ѡ���)̊8��LK@��>���a�=�'�P��>�7}z�t��}����Q���?��|a������H�Y5�Kiv�QkrP���Bz�E�LI�[��H���<��D�nSNB�Uy:�n�f�$j���@��x�#�Tݞ3�u[����\���@��3��L\)U5�b���
�����A=�>�Z�٦ZU�2�&�����h���]9Ƃ�)
8]E�����?�gazPD:���l�'��C�
u�u�-��>�:���F������Q�wyg���Rx�i[HgG��kӫ�kݞ,T[O􆍮9��ϛ��Hچ�8<�8���t�͢����j��������Y@��r2�(���+�
*IP ��/M!@D�.�����'B��I�g�����d�XVf�Xl
8&���v�!�͔��G)h��JHLV	C�{Ј~���z��7ޡ���D�t�"�� ��k	�����]հP�u8[D�UVgX��c2����X_�*��q2�S����ã���8����Mz��F)4׍��1E����gd��D��榜`a�W����'xyA[+���ٽq3��!�#5V�^S\�d\v�������;lw��+�|;EQb���	d5�Ӄ��H\���Q�r�-D�+��[� ��L����d,���x��=`�bn�8�����xF6bo�������#4aZ�j�q������\b�d�� lf[럺#;�e�yp¢� ��@�P��w�i��5��bf���.-9�{W�iJ��X(���%�!dR��A���e٘_���G���m��M��b��P��)m��Y��%C
��@1�������AM��	ê��
�W��V\/: �dL�㈙;�rƸ2~���x�z�\�Lt���JC��#����E�&]���@s���7�&�p�_��Z�Zݗs��0��"g�䟆p������c d �䠾�Yn��73�$�v�}�d�	�	���{ဍ�˂�bj;Ѹ��yil�̫�?K#z������T�5��i�̀�,uh��������OJn�]���Amq8��S�A5k�z�9}/��A�t�0
vj���jp0�X���Ц9>�K�%sU|�$�/�1��;��d�ʛo�s������.^[����7��R3$�����{��h�c�0��=�z�	���>ȟ|��2=�yx�H�-:�4�f���I�b�N&�P/\S?���(&f����u:eC��n=�jHݟ#M��������Y@��Y�Vȹ��`u۲(Y6�M�X���r���e����y��}��ť�fZ/�b¥�9�*�R�y�Z��}w�������Nɞ&T�	��m���� O�Z�vݧSd�}(�s�{�t�e)a<�h�壀�8�k>�tN$��^@��ж8f�% ;������	`�L6�i!���9�q����ڙ�;���Z�XƷ>�-��ޔRO&#P� �����'#>�v���.��e��}/^�G�$��h4|�_R!\"��}+�_�|)��˷T��Ɣ`�s�_X�ǁ��D���	0/=Ml3���&�\t�� $�,G!�t��C~͆�3D�v��Mý����j�ľ�-�G�k`��L��+�+�vڻ�E]�,()^��6}��kR���f{�&�Դ!C��ʚZB�.���R�J�WO���M��a"0+o����N�w��#p��$g���B~A79�D�bE
�\l3�*bO&������g�­PP�*��M�M�o�X���?g]՟�Aw��;�]g��W��E�:{������py5�|��em7���=
2�=����}v6ض��8F�iZ��D��H�f�L�W�%�_0 �8��[�_��]��Ϲ���e�O䩵�lWuNsU���c�կ �  
�c����K�-kl�!'ZT����D���w���x�"�J������2QlǡN�r=�(�3�ue8�m�@)���+�df��L�3�/Ñi�������1S���߶����eվGƮ&��<�@->�\��bu�o�'O��N��}\.ݏ��A��\�����J���e�=�­?�R��S@��H�~Lk�LG�t+hzsf�9�xg�Ehk��[��	5]��xk�CXE�j�v��'���oP1"et����]I:��0��֭���c�����%��^$v~̆4G�S���xC���%ѵ��"��uU�1�ߤ%'�4d�tg��,��l���A�!u�2�5'=ɢ)u��(�ʱ����8#�?q��>!C������P�z!^:��mAzwQ�/���������^��x&J���s$Ѡ�k:,=~�����6ۓ]7�!�H�#> ��������y,�z
H�RMN]U�Z���{���y���6|5a^\_�QO ������h� �E�OxB,������t�/�`���i��nV���G,	04��t/Ip̂���%^]D��:��
�5����)Q�r{Du i#y"y�_�S��_<9���9�Dw��
-��D�v%������mݓP(�A6����.�T�I��h1]��N��|����qQ}� o>�ʹ��9]��A�'�/�~��}0��55I9W`��n�	�. �v�mW�����Zډ*XP:%��P����^�AO��,�`��e�$/���Y�^�y���n>�xZy_[�$r1�fj��Zأ�[�����b%@���`�K.�� �q���'���30Ȳ�#?��>�@O�8�̩o7��/a +��������Pۙ�֔Q���S����������6�X_H�KX/��L��及�hos*XRBs�{{������^Lˋj5� ��yd�7
E8HT>?���3��`�
��Q�w(7�Pu�� �9�y�K�:�++�?���"��c��a����d+o�ڷ4����,np� 搗C�^�}��'6NF�y�Y��:niM�tfz�X�T@x�.j���^��F���Awv ���6�1�ڿЭJ�2(b�Af�b�%�:/��6g��O+!�J�����0u�~���0���`��[i1�a"䀤�6;�	����PG��l�Z��b'����f�`{"L�|�Y0�����G�WI��Q�\�:s�y��	>���.w��RNBe6�#ԇ5f-�ϣZ�i�T� L���m4
p����%ô����q���`����t�bP��zY������Z�c]Yi45-E �)��86;��T�]��QҼ_{�aw�h�����a2��S=@y%�=�� P��bՂ©�'�����SJ����Q���A#��<�&�}¬�Vj��[׾����
B���1x�A�u�N�Y�?ձ��a�%���LŶY�[)&�A���=*3���U�q�ݑ� R�"���.���ܵ�rv��?�a~�P!2��)�y��v��^y�p9��mr��|��dL���j�ƑL�a郮@A��byDm"�% ��ͣ*��B(�y ��ܡ�*���K1{��}�m���� ��3T�k��S�52����9i�Np����6����nÓ�I��~� �{��j�2�������،�����/����wD_��ҡ��~x�KI۵�/��NC�J�=Ҿm��!���>�c��]˦}D ���Fw,ʁ���ZŮ�x.�(_Bx岵}����i���́ߍO/�毉�~&�Zp�fJ�,�v!�x�t��`�N�Gk	�� �l�fy�#���C�����VrW�Dq���΢�3��)�3��gt�t������ ��,����7���Nr��zr�l/�%G����� �PhdK$�+�K�	;� ^��(.˴8>�aX��3�����r:�1b�m�X��T�����0� �)�_�e�q��[I��Ml�>ׅ��Ì({��u���ﶱ�=�s�)W�"��I� �uQ��	6���%0���������|���k�h6���%���נ��M��Zc��h��P3��g �A�E�EV@��=��¹��g�C�^ֿ:â�Se���^X��������f�#-/�����r>l�b�1����hK���ӿ��Ω�"2N";�����\��C=[\{�rU��>��}W�Z�K���[��E���TS�G�,~�n����`�ꈅk2,��B�!9�&2�����V
����l��cH?j})S��;������-x��䪌HWv@�h�]��Vڒ^~$?�T��Z�������j��!��k�o�Bb\
�#�Ն,��O�ȥ͡���'p�s+�Os���ٹ�,���������,�C�D�c?G�w�D���w�]Z�{��?�ާ����}�|'�ͫ����!k�[�*����I�ku�M!����J��-�Gܑ�k�C���&�x����s���e�{�oo/&�ސ��əQ�at� ��?,\L��h8�c��cؤ�����ݽw��=-�����N|��X�|k����Aݩ!��r��;+��k0�DJd�����餦��w�M�5�}���k�9������I����~�;����'Å��X	&�/5Ǉ
����:#��#��MP��^iP��~�t���H}�T�K��-�|X5�������H�A�����A��m3ש,��`.�W_����&k�|�=q!)�L2����t�yXLʄE��F�j�[Q���U�X�ˎ�o�I�O�N�uG\{��N���vr��9���nB��Z~\nwk��n|alH��i�]6�7>.T/)
`2s� ������
��õ�� %��Y�q�ȤD�
l.D�bK/������Zy�b�ȋ-�d;,U���Pfl��C��i��lo/a��=u���;�<�b������v��E�i,wn�M��W7�hyq2O������܂p�N��1>��O݌6?�ly����6L����:����v���9��ܙLϖ��`V���s�@����9��}庛?7�(�]�L�)粫����{��n�?�wX���j��*�1���	Rӊ�h�xi)�,t"�'���� `ὸų�^?<ld|�I�P:x	���*I����߱�1���J��jI�0�G�ʊȧ���&F�����t�֑S��KB'���D�;D�\�b��<����ɺ��hڣO��D̨v�2`�$9���eI*`:�y��J�<)�okb�gl�?�Eh�t:�����i���TQ��Uln��HXȁ����B�Y]��t��X��˾�U�Q��K +���X ��L'�v47�vn�PI�Qw��r�RU<��EB.t,k��YT"��Q�d^r�3�Q`����|g�	��?�4�q����p��ɍ����d��X5��%����B"s���-������ֲ�έF�\�[��1Pm(f�W�����ֳôԭz4�n����r�?�Wl�`�Nu�# ���nEp��SHE'�Y��>�2.�#yLr���FZ;���B�0�3���P����b6{��-�}0�G>W�a�Q6����~nd�5�M7��|��~���L�:!�ɇG�|U6ג�e:G7ClQ��n�|X���������}���߬$DGc6�n���4���%y^�����B'�];-��,"� ��k��9���q������~��w����#ڢs��=v��n�5v"�k�uI\�=��P����c�_2d=�(n���`��w�߹�]�wb����Þ�Z1����#�b�ikk����.0�w)*W�s�r�����K���+"�h�X�"H�&�����
?9���4�#� �DK;;Ew������-�{I�J`��1q{���_mi+�V;(��"���׉W�L��G�@uӫ��B���U���p뜺��DxP�IHed-��L���J�N��; ����d�V s Uh�Sߝ;i8��ġ'�.c)4vM�U&W+�bׂ�/���`���X�o=��(ˠ�RYrS�V$�z���ab=F�ٳ�(Vx�.��e���RzT\�+c�gֆnӿa ���fLa���TCݎ�O�x~g㒹��G��4$�+M�$�2'��!U�Z�ww_9n|�a�QhP�j?�1��:����lݒTv�#p8ò��mmb�[ɴ�͙� Z�k�!��%��b�MyT�.�g�rοx�,X�4��){��o(S��9JA֠b���#>��-�",�15z �ʸ�/��8-	XR�����`2+��ľi�y�Ѿ	��
,zX��rעq����[R��/������BN�ٗC9܃G�
i�p�rlE�T,��ٝ�?ē����j���Xw�K��x�b���o]��/���e��'�d�&tT+H#�ó����2t��*֥�px�
�n{@v ]�Uʃf�A�W��J�c���a��X�*��W��w@/�iC�(��m��UYٟV���"3=���t�shgp�&$Z���7C�{�M�R�V�Xk�����Ԩ\�K+��O����o��ٮ�K �ʁ������K���������ڼe�8�=58�v>lN�� ������4�bQ_����7��Em�<Yj�m^��+ �n@�^3ܸȒ
��{w��B���������D�>( R�Cl9Q�;eg�G�9�9��4��B�rĵN��"i>���\�/ �7��eq�=y����k�c+(/CE�u/;�|��~��d�E7M3I��h�4jD7�HR�l�XT�����3�v��󚊶�fܽ_I�覣�(�! m����@��B�}���#I��� Z$`_���!2��IwƌM����L�_�=�6���+�!-�E�݆�Je���?���Қǃ~yf(�.�|-$�Վ��'�U��p.���݀�����qрES�����:k0�'��)�Rx&͏nu�u#��34e��/C6�14�ݠ�����JlU��&!&���������7D=j>Hx�W
����D�n��(2�	�H����,*;yk��̓.�+�^e&�6m�&��t��l��x�bGtk��:�0���:�<v��Pm�g�/x�����0��q�L��᭬3�m��}�v]?ܠ��~Gg�L)�`����!����#�dֲ\�%FUĖk��c�<���4�HO�2��zr, ���eT����5�c	)"��L������<�9�{t�X�1^����#OiǇ�� @X���8�ў���j�,�����\Xf��+{�8�Ł8aɫu<�9��^��h�.1�T�}�D����R�h�o�X��[W�S��&r++�Cƕ�sJZ9����?[~=���N�GlS�'�Q�p ��,�G@�p���鯅�C�w�������J��W��9$H��K�7����TnU�#����&<��1 W��L"�~!��@�م��{�|��׿��1�-L̼e��(��otP�h�Z�W����w�28Xsc/�|V;t�{�I�f����*����s�ub^�S��3;�;� /�ۿi�j��oǂ�@oQ�}C!V���D-t\J-9�,���m&�&zG��P`�����%d��j;�e��C/Q\ѼK��xS����
�������2e�ݬ1�n���feq� ��d�& ���E��|_G�.��g�`�|�����l~�7�2�Ô�[��#�� ��5	����� As��e[��>(X�ꄿ�K,
4k�Y8�-tjqaS��Օ��?ܗ����w��Cw�aү�Y�xV4ڼ�b$zy��4�����W��aP;y��̳)�|=����D�\��Fsx74��ՍA�)2K+˱-h��S�I����!�a���\����W��'ܷ����|�5A���کy�I4�W�o��G�up�RX�C���B��
�u��7����]DI�Q=oϐ��-���֤����j��+t�Ke�?�v��3�X���3��w���� �Ժ�dB`��5�k؟���_�!���Z/��.�a|9�@9� ���u�!�-3ϯ�˄]���ڽ���&���Q)��h%|r�Jd�5�g7�l�����<_�����l=��E]�6t�Fs�u�n������;)9]����sH�9����@�q��@�����t:=ϝ�Kz�]�j k���@+}�/��	�53,i�Ī������A.I��ģcP4�i�g+`���3�s����a�9�\�b�����#%�{Ԙ��QVN
�}����:s�)�Y[�^���H����6xm.�6��ܕ��B&�2�'��٩���Ò�_�h>0���5�h� D{�V9
UEo6`e�
�#a�R�{[���'��}wz	h�v��Q���5x�^�5 B�#�G�F$m�J �f��z<�ݣ"���;��P2�ѝ� =��k�m�´�}>B������u0�Dǧ�G��^s��dф�K���?�-(*LW���5��wV-j*�"��Ot���]�����6��j?MN�C%�����1�l�>�ޑT��S,s�C�9�63�~�����*T�lq�y���|���)�F�A�3�ٸ�n�I���!�!y�z�3�7�ߔY�F)��[��kF�U+^��e,f���%F��x�"�ԗ���(`�^��$+�(b.��f��$�!��/(㐖0|�嵕Ύc/4Dd�b�KG��d^�j`�/���xAnnE���S�� ����9��%$Cv�f�z9�	���́'*dS��ӝ��Z'6|��X���4rͳ0�[m��zD 2�OS����
L�s�`T����I�xl��C��"H�])SR2x��xIm��1���tJ��Qn�Ur��B��h�{W��**��2�p2.��eC9Zy���|=���kY��);b��č��=����>i�!RD�>��A�)Yt�<{�@M�ԍ���8&���o6��fE7^����h���PTh/�\h�9�N�v�VOO�в+��(��M��4�PA���tJw�.>�C�=�T����'I�]�7�#ݖl'M�8�?o/`m����Q2��8J��$��v	+�4��[H�rg��E8Fp~���%1l����K�=~'e��	RL�����k��y&�1����ݤ�]�++�=[b�N �7O����͢����U��f��VH8,���M*�;�o�����Dەhp*t_(��<�[��L��v�7�ս�e�H�*N�X�3�i�x1)�P�rcMq����͘bE��U����=8K�o8�\�D`�/��<�v���L�\5�y0�)����g�f���}*��0.�����b�|�\t�͝�ӉOk��ۥ�Ue�!L��8�Q�81��%�>�l��qYC�u8f`R����!���E�=4���4f�_`*h���zb����@�U��_^ȣ�H�D��a��c��I�9�d�=S��R��*'�[K���ȼcm!`�ۡ�ڙ�����{e��>v$ VdލRT�+�Y&���b�H�ԅ�Su��['x$���G��F$bi���&+��?���r`P���?GK��7=��O�L`cܷ�@���%�ܤ�!S��o-^�O.��0^��co���g7 ����?8��� g����ތzK�ӂ7�:�XP��["-u���%~�ќPA��0�ܨ�'B�V� f-��Z@@1;޻^���oAۃ����v���8%/C��z��U@
]uz�['�@�j�����\;����Sv��"`�l "��p�Ŕ� ߖ]��h��h��,Lg��V�o��D�!�H�F�(��^�����sĺn1��2����"R��w�F�X8i��f�
�
�Q�AP{���%@�ݜl���um@}�����k�g�G�1��V��e��tc�<DI��5Z�#�JE;�m�$��P,*ҩt��b+U���z8�����E,:kRQ�_��<��i��"��Z����[Ɲ���,�{��C
�>�sp50gn�K�D;~�	��������yW^�
 ��ÊʍC����n�If�@綨�_���vѵZ��zu��5�
^��u��Y�&oO������|6v�|�|����`�X2)�~���[�x��ߴ�2t��y�V�sa�Ѿ��?�/��4��Hl����zpp-�maU~R\
�v:�n������a�J��a�0�)��������8����E��iF��)E� û���������`��n������O2�(�c+�#O�o�:o֫��?A���>)s
��Y �1ُFU8��A��xd�c�s�G?U��d%UvG8��ֽ�%_�L�>U��YH����w�-�/�m�"�����'Ak̠]��1��tٜa�ْ�jED���^�u����H���f4ے^�����	�ϫ5V|xǌ䮰
VS����+��R��q�W����������h�9��8`H���fT]��M�M�����X4��K��}�C�^���U0M�%��n��`;b[W^Oܴ���j�@�.��F��8!��@��
�Ϯj�S+?F9�g_9�-�K��.v�c�r���y�B!��$v�+Z��Sa�(s�1�� #�������T>4|?v�BɲX��	�"��3���W���v��gqFH\2��bS�/:���{��Q�T[�n �Y䂓��c*]!�^*=�r=9p���~o��w;�rB��%WB$���N���7Wm87�A�P�ҍ�zP3��y��*'DIM�(�O&̞p�}��.����;�0k�c=�;�>�LiEP])?�S�{�0�Fw5��b�ƢFÂ�P�0SB2�Ǵ��z���I��	� @n�FFN�ș�0؏˔��k�z����}�ᢦ�C �1}�' �C�!��|ށ��Ū"'�PmH�U���P�P8Y4���A�#SJw��3��
E�*�)pC*;�8��.0��%5(s�#S���[�p\�*v�۴ �cY��þ4�r��Yt^n�A8
p�	��*�j�sn4�l�u8�h�4W�M�a�f��;�'�Y&D�8`�6ͫ�?�Z��{Dq8��T=r �)�i�s|��|7�2`��z��z#�6�>��̒A7���-FԨlK�:F/��U����T$0�7*��q�Put}�a�}'��f��ګ��B��cXa��;*�q,`ԥ˗�ẸC����α�7�!P�c������=|��H2UJY$��ŘnE+n���Q��>�{u)�k�V�b�,���m���o2!�m3�S�\Ȫ��&��{f#�r��� �h���&$B
�.hWE��Hz
���{̧��WT�,]n�\TD/�"#;7v��b�o6�W�~V���M����E�W;"Qu8.�V<�pWX�_'H��"1�s-�`�9v�D���[����xh^+I�ß?�c�T,�@D"	�������	k�H}�b�W�~�8L�U�tq��|l/��e�U�D*xlA:��r�n-ͨV u�W�����y���*�;][_p� v��S��^y*��\a��Ѻ~���_d� �'6�9F%���S�|:�S���/���A�%�~��7�o�e�AP���[d��7�%�����h}�CH@��k_�����<�Bi��XU��k2�� �}�m��?����A���;7#ܤ>.9��%�NcL�75���2���4�,�_�qs1c�*r@�J��	�#`�6�FP3	-��G;�4�q���7e̔6�g��І�Dy�g���a.�DSG���>�w�C���=��S
�g���;ț�p�M�9��C�wݢ����i�i{V���ý�k����ؐ c�ޕW'�j��Qn��S���cJ��F;z���<�b5����윞s/�a�
DtP�#�arh'�j'��S\��:�1?z%u*`����%��Q��=>4b�k���:��>�z5op�Ѷ(6%�@��y�Є&�l"IO�^�pls�݄��#�.Ć;���,u�7C�o��^��ņ]��9�	�_O�c������d�we�$���_� ׮&�m	�Z*��Ïgut �	�rA�f+&0�Y�L{��GPwG.û�R�Tb�v�4���X?��e�p��ua��y�֌k�f<�ˁ(vOJ��w*�@`�C|3#{��O����פ�,}�g���S��&]g�R�@����\���V%(�Qә���|2�o���_U��.�6O'Cq�ȭ��x`#�z��M���u����:yfD�L�7���iT9&F�R0��IH��?Ie#f��O��k��.�)9:�|�w�	w����&���f���A��A�
M�O�8ZI�k+[��*?�P��9p�*��b��GB��`�-7��UɉK�Y�C\����]{EC�R8hF�+*b	����ah�A��AW�tl*����Q���nDb���4k����&�Irn�������- �����1�BEmj�X�se]��]Z���`Dؤ��dS�KK#�k�랠Sw�F~�|���˝��aCHQؾ\��O���[�T�N�'<��ھΧ�r��1~F��PnA�j̲�is`q+e�Q�Z�@����ɗC�Y2}��!R5n� q�Bd��f��}��t@	�?�o�W�z�β��e���rN��S|�?75��ߒ�u�C	Z7�?�hN1�j�A �("����B/K���Ʊ'4���ډ��(h^8������q����DR���d�8�b��Y����V�ÿf�\�g��l�3��n�a_M������Uu�{硧�o5���.��+�[w�sS�z�z?:g[� �c.�l��k�g���[��A8y��!��pB:�򡣉�t����+��CO�q��[q�ۑz6A](\-�T&zY/1�)wK�x�4���������;��eʌ�׈7G���)p}uhQZ�p�IE�Y�E�{�����M.5R
�|� ��������MZ�F>�m�ι�_M,N/�]��!�o�ܛq�F �;�Y�~��ԓ�(������{<�1S�Z�7o�O�"[P�%l	��	}�Y�V����M�� ����r���ߢi�9QG� ˾���F'T�6b�����x���^��	��"YYD�k��>ֽ��\�Xy}��{f�����p�/0���z��������al�)��9!Ұ�U��	<=/�ɧ0����s z�����F,Te�w�%N�;��^x�}�Ȋ�y�%?�(�-rFk�`�TCQeq��5^'*��E���W�Z!�n�ʻO7���F&L��0�En#'��_��4�O٣xe���A�����N�uE��rx���c���{����A�MLR�.#����xצ���J�$��`J[ �V8�5�K������GE���'�#W��oޙ'�xrYyO��5$TV+�E���W�����.�c��e8|��-�Pp9�)߂�f��8��cMbk�`X�as��0f��a����oo�RV ���DI��<�g!MU�@��қ&�6i�������,�D��U�mL�t�i��*a�Y�tZ܊L�z��$�/_�r�_��X�,
��o+8#�	 �kF�'�ܾ�+�`�\ ..����2��1�N��l�a���rH��潔_Z#�a+O�'���W�x���$\���;���
��M�l��sn��B{%(�EƷt�����5E^��;�3d�0q�{�	=��كCh��L��}���p�>
uwvy�+g�E���~���/�C���N^(��{k����0Z2,}A��s���EN��	!��Y_Ra{���AL��h������%������8�~򳃐��e�rx�����	�s�!v�E�	����]��G�Ek,�Mk��:rr�A�M7��@��&�~�����:�a�+G�c�ng3�7��K�3d���� Q ��UV�t:�I���M`�.B��9K��|�������I��e��"�Ԭ����O����a+k�����b��;�.y
�NX�R�
�5�/��FT��c_U����͖2�%�_�z�|={5���_��K���R�tM�*��p�V�N�x(dy�Y�gJ1��(l,�� ��$8�u;H��p6�5�0T0$�3���p�s8+�0l݁�\�cA����L����X���q�+ ���γpa@��zd�0���=��A���+�j��^2���+D���<֖�8�_֢ê>|Pӵ
�I�zOCx�2�A���cM���Y;�D�	���YB}랮ft��tӸ<��S�lZ�\[�wy�Lw!��՟3=��1D'�G���C�H5��O��H�vr����t�a��W��.��{^�)�T>tSn�Ӑh���et
�#�Փ8�g0B�o�ک�,�g�����/���]�p�٘o��8�E)��(Z��ՙ1itoo՞E���D�p3�cWi�5X��q�q���Gބ;Eq���6���̶�x&3�*��Y	�d�IzR)r�j�H9����b���A8��'��[�^���珁���\4�n<Z�ֿ^�B`��7�1k�����LXF����$�vE1�ƿ��k�g0:~��=�6\n�\k��A%�b��Ι�F\�K�G��d���v�6Z�e�T�a��-�0��lq����~C�l2)�*@��U��B������B�EP�1#��@Z+�K���)��$�=�� ?b��y�w���xh�����C��L�'�_6=B���>�(��Ǝ�$T=o�UR���y$��١�`P�ޟy�N��fPET���A!1�7�xm، �8��	<�a)b��o�ŵ�?��u�bmo��:�*��h�}�y�����wh��J���,�~�YD2���g�@�����M�e��Y�e���$E����f�AO]�s�;���̸�`L��8���5�`??Sz��t#�h\���-{�+K?"1���=�4�%�${�_��)U����h�,sK����b�37	N�m��I$C�zdu�9l͑�5��B���9@Θ^K���[{�ǃ�H��䨒�V�G���Xi8�7+Lߢ1-�͆���ô�<���M!z��E��&���8�j�>~FE~�x�k��qx�E2-�%�-54�4}���g'?���e�IA�bA�v�A<��R{s,>rS�P��7$h���@&�r�΋s�_�i" -ٕY�eR����
�F��*��#j�1z���o��Ɛ%�~L�
�?��Ѿ"��A�.����4��ʊ#ٜ�@"��Y��`�7_](kMP/D�{&����s�.$���q���Fn%u�!)9��[1��4ٞ�������E��60�k���"���� ��(n&�	�A���&Ŷ���O�35'��~d��Z��鷡�Oj�b��,v�8���v��)��Fe�6%�u���Wl5����,��ū���7%~�	'_V� ����grN�V�x;�
Aiz���[�o�����hB�ܭw��_�|�O���h����f��ĵG��d��(r��w���x{tbz��O?�}���@���J��x"�*��iEX���U�vq���ߎ�ːI�=#r��QKQ���i��K�DH�]��P�/.���OB�Zt�_!_�P8�$B~=a8c3����`x��)�tZ������Ν��vh�{�,q-d��q̑%� T���g**%^��f���*N	���܀P�.���@j��
�WJ̀��A��Kt�2��#XI+eڵs�����d��q!ڽ�ќS<����q��]���Aвex�+�Km��T=�N��l��;l V���6.�I�o�7�r�5�`V���Ű��Lw�L7���c�Tլ����g�����uT�3�����B�\��/�ތ��'�f�O�n9h��u���+����P���D�d��%Ԃ����pɦ3�Χ.�v����5gŢ{�l�k�X�:.i׫��;l�:㒍,�����NZ���S@.-}t��ï�R;����a�gM
9�0��C�Z)���K����CK�U�*|��$����|@(��¹S8A]�~�����Pɷ*��#�j�o��͹>�w��
j�(�r߁�0J����K����yh�v]'��@�����?��p*�/ڔָm#�׵hC�#����8N�x��Y��W��������eJ�"�3N/�kCg���D�jQ=�����g]����Z�5�ѥ�M4E��3J�KK=-��_ �_�o�i�E?BP?�b�|'W2�� xK�-~�YNDV����v����k�T�A�l�:�'��g_v��a�V_�}�f@�.֧���׃���4�$��#�~�^
�uـW�o�8�N@T�[/�����E�Wt{�c��� ���2-��F�֐2���Z�������s(��aq_�N>3�F��>��s���m�`�gr�;�E>�S5&e�Es,���8~��HZ�w��-�5M��}$N���9w�A��t���=.>�CZW3��۴99}Cx��6���ԒP��幊���0�;�/��
4��o���H�H�d��Eӕkqׂ82��T�iH$^x��K���8�ߧ�9jX�51��`��ɻZ��2�+Z}lS,YnpA�����G,!P�������c��(�eg�s�h����ą�Y�|���S]��V�[����MI�5�dU��BJ�:>jL���y��jݼM�r?��c^9��R}\��bR�=�Y����v�UZ�ِ����ϴ�<�2PE�`������H�)=��,��E<��gla��Y���fh������d��e���T�"�G��pI�I�{����_w#5����pAnS�4�����K�c޼v�5�s������Z��K��w�a���u�V�k�k
̑T.��M�%`}Q�\��P�񙃌ٗL-��u	V�<EO"��ɬ�3��]U:�VW��(#c�ܚ����p�Ş�q����W������ӧ�E$�\����e��D
�i_�4gro�kɪ݉o��I�T��a`�ц�F���H᲌�| %����^3�ĺ��пfE0��C��Q�X��"f��X��\FI�V%y����;�4��U�f�� �n�`�_�;�.BP����[��$G��N8(f-D#q"�h6����idN]���U�&�`a��a��@((���ʰ,v&6b�	%�ټK/0�!�1�P��P����a��b�V�oJ���2�7���#
]��J�j��5�f�/���3�&��C)����U�bU��H���~���p����/w7V��ks�2p�����E;��a3�R{��:�>�X~y�����F��SU\p��4x���"�0�7��''���P.�3�|�+��B���b���y�"�G�(-&�_���$�g*�/�9�`�Yы��f[݂�N�ɦ���]/�e8����I;?��'Am��1����֥�HEp}Q���<8��eONk�4{�}
��g�f��2jP�xy00&��m��Ef��i�U����rje�:�i|�%$p�+�ٓo� �m�N�������Og�?�^�g������h\G���NFb��gb��h��^p���Zɽ��s��I6�<ޔo
;�Y��+j�_9sc	�B�Xr�[p�h1���aN��)!j-c���+�Ad��FbuTƫG	7�`������&83q�~\�j̙�-����­�X���86w��ՎϬ����jO�WH'	��*�/O�V�7Q`�p̦~M4��Y�������y{�E�z���`Jb��Z���D����fn�g�$�2��������{W+�:���]�rf�nJsB�� d	,V�-�(I�h,�����krƺjMe�T4�c��E�i��Y�jj V6�A=�˖��m3l����;g��#��g�V����R��в
��I�Rz�9�,+�=�S�(tp�б�-�ЅT.FS��uBU��:K�\,o�j��I	���*�	'����.d��>�G�\�}np��z���m1ڴhyCn��Z���T;%�&�a��� k����Y͈�Ls@������o����U
 �{���9�>>���m�G"��Fq�}�u���T��tM6l-`N��FA'�J�4��SmzM���|E֎}a�CBy�KO�A|s�n �5���n{M6��^p�L�E\�����qC���;{�c�b�#���r��X�G�C��־Π.����6����Y��P���jT{D��d8i������4��7��9>�ݚ3�G��P~8�v����8V=U��"����b�����.5����l}� kS��;���~[���;3)U5������V!8M�&頋T����X��I?�yذ��2*D�^�+)3U�G����vL��J/>�~M��K���Xa+�K^�V����2Ps^|>Ů蟯q
&��5s25'N��\��J�<x���P0i�$��3i66U��ܽ�~)md�Ūi�r�Hw�M�9�-s��Fq�g:E������o���㊴�T�[]n'L���l���ǠK�D5� Q��pٞ��Yy9wO�<T��ޜ_ɾTj_��?sI8���D]���t�{ۉ�b폨P��s�-���x]�OO�)������;1��҇&���p���o�����
�{� ��sCh(4�8���r#���|H����^G�]�����p�k�R��8>g��"D�C�%X��Q+��K�����F�[<�Ƶ�N{�Bxfջ��ܜP�<
&�d��N�J]���hEbT����>B�1�Ű�eҵ�_IoMrx�#Σ^k�(�y��YPƅ��LO�+�~8���+�KVΙj���r�+���X;�)Gl�������x�2�#L	�з-�e�Xz�N���3bl]��ʝ��A���O/�����%�z��P��煚b�|R�ܯ}<��
�%?"�E5J�չ��5��% EQ�\�)��(�J�["zsj����ox�16�D�'��{��:b�RV3�n��0QYT�i���	�!l��:V���Gâ]�ժ�d�(���_���`j�ѵ�� 5��ϝQ��x	`�Q:��5�A`]h���ӵW�"�3q/��ET���rҨat��`�Y�;�ҙi�"i���NV��~ @�H Ye�lv d�[�ӹ��'!&B׋K�v�0%�͞"n׃eL?7TT�Ɵ)Y��/����z��xG��.��1S���ظ O>�r���wF�
G����y�}�䙥���J,�^��\ǘ�I��~8���~<���D\�GL�a6�*�
iS�D��{�������,Ml@�aHz�2s��qp�C�G}�/��`t�r���p
ns8��f�P�W��D�lC~`BkSc.6�
lghu����1�w[eM�%��B���#k����/ʞ�{��6��&{���m���.'q�)ߕ|��j��a�1K�m�k ���֌��)j_��:��`1����j�jń�LiLR'Y�- \p	V$l�Z�Tyj�~��m��h}48�٨��@-�/��� �_�.�[ �I�|C]G.y��e���?����_�{09��6�]R��-O�/�C)�D�;�G�����#j?ۂ;����u	u\(����6;f�e_��h`K�\�H�jC^�S��Fg�+�k��ث���2�S��P�%e/`c�h4)�cGP`�`~�^X��ق�4uQ��{��7qPL�'���?.��L^U�o��_��\)�[�TC��j&���м#;����E�R7o.�d���Uq�Bь ��[�'��a����cf�/��gB�-I��+r`���5Ϗ��bA'����*��pl�CY�U�ʜ;	��A{%1��?b������;�ҍe��*f��.U��D�����&�+dt\
�*�Yо�������BdƆ(�G�O룒�Ծ�����U>�Ч��>���[9h�4D��Ωo|DQ�X�g����|h���Ï=?�q���=跒'�������O�N�ʏ��Q�c�[⤵8�Z�Ss\�J�p���N��N���nE��)} b�"�B!���>H|���� ��<�t)+��vQ�`)1���'�ҩ�C|��Ѵ��iPi��مs���=�הq9V���P�<I���E q�%�n��u�i�u8<H�;�M�G~JS�} �������L8 e��3bI
_6��n�ɩ�2�u�`�
B&R2T�\�/z��ۗ��c���?Z�[�U��?�NS^�p����e�Er�-dKg��ȹ?�	�i�l�,Ğ#�"Vpd'�؜a�� �HT�n4��ǳ ���bU��A�BS�����,��Hkp�hi) #�ї_z����.��X���q�t��Q �Yz���zћ�ƃ����p����.c���r�b~�6g�yd˙
�RM�s��ʪ�eݥ/(��`z�o���g%�[�Vۻ��(�tLڥ������^\r�8ꄽ�2�ۅ(C�6�a�=�No��7w��VJǧͲ��h�wx�u���2���([�����7�9g.j�T���<��H�?��>rs��x@_�3�B1�Tr��; "����}jQ��.�;^�#)��Uen����;�\�ɛ�����J�y�W�ێy���ԵEI?�1�4$n�/^ms��Jqf>d�#�]����m':�w
���F�?���B�����̞��{�LE�:����2�8��7�~�3L=v�RXc0����(c�s�%f�B��v����r�/�V��*o痚��!�c���5mLzc[^tD�KȌ1C�	��b�G���~�5���H�8äw�+D�4���7UW�{q",�צk�݁��O�UJ�O�	|%��Z>�"�x��&���f7>�QA�AqbvGj���jT�w8{�-G��� oF��K5��+,�8��f^�c�0�z�:�1ʧ�aڟS��;=��}��T�}��L�m'�q]���d�]FI!����r�$�*
�.���DT?]crwP�F�!|��z�i�\��5���ee���R�v:qEE:GU���4 ���^��?z;��b��Z���Vg�g���x�\
,I�����Ej$����#k:�m�4�W�D��&|e�1���9����]u��7�wĺݣ�}Q����<��;�!��M������B/o�M��)��`Œu�3�$�;_��D2�AF8�A�OG�#���k,%����?^]����c"O���Mr�{(�Kce$x��-z�=6Zk*,7Z(�[�����&�f�'B��M����%����*u>���T���`tu��FkЏr%�1�����F���k����0����sb��c��H����}�+N��"��P�~�
Q�>��7E���Ԅ��7EE��?C���3���O�%vo���=�u��>7:�������M=��(�m����?��G-�ܓ����H�Ì��uY�����i��	x��Ӏ�꼡�z���<�?i����u���=�ٍ�8�=}�� �pdh�9�"��"Vq���:j���4�ѭ)����݆�as5]�k޷�~�\��l��ܽ����u�$��1��.��:K�{Ǻ�2~�`�Gy,&�����1|�'���Ǩ|��^!<;�wR�Em)������}@(�sތ�3
]�h��*F�Hz��rgΞ��o��l�NN��sUe,Cj�*�@�N����g��n���^�q�q׸N�1���凃$�����NW��q��y"��U�b�ۍ���>��]�rR	�r��wo��|�"(�*}��nO ���]cg7ת�[>�촂���=�����d�H�T�#�d�}��1����#��&��D��e�T3��{��/s��[/IRv�^jՊ1���g��Y��d^_��5�:�O�8B��za�{��N���VaDP�ɝ&uiJłF��A�<�P��!���~��/'�eS�	�l���v6"D4�BR�	]�0@]S�a)۟�F��[��S�L�9y��N��ΐ�dH�4D S�JDf���)Wسɉ6��PaQbȧȾ�ȝ�� O�����:�����N����̨*&����fzB3ڹ�K%|_]3��`�Q��æ<752�� �#��������H�;�����ҵUS@6RF]~�ٶ̘���2����Q����,�.���h�!�G!��%6Q������GI�`���i�H��m���6e�d�?.��D�My�$�&��T��	�bL�m�:�RG�R�͏��
s�W�vN�VL�sy�RL�b��B�b+���O�ق�I&z+BWR��Q�*�.����!7w�c��0F��)=���8��,$9i|S�J;T�	2��kp�����)Q˰�A3��_�kzfW�F
�v����J���(����+Gx���V�.�^CP�x͈��AK�O�<.����T��$$��6��=���h4ch
lһ������'B[)�\Owk��� �x(pYs2�H��rI^0pd�M-*�7'�.�|@R�ρ����Z���Qv�P�֖�끂H�Jk��{T[���;���b&g�SE��g��Qِ���J.�����3J�2��f����p�hV~F�֤ bT�.Ѡo�4eS���5R (��ì�5,�F�!M��RD����2���㼖yqa�<a�<�⬥���H;&�5`�2J|�ɻİ3��\�߀�ǡ�&(�
����?��\Es'��|.}֐��(�nA��.ݟ����\h�	�7�����ܽ���Q2�����U>���J5���5֧�dwFH��~��b?��O�Qy��S��>G.�T�v�����\��]*��f;[�����=��ϑAFL�� +Z��v������^�L�YA�}�������L�U�>sb��a²�<f\nW,y��:�㈒���qd��T����_�츘�1AI$�ļ��H�")�ǤŨ�5�:�u<�2:cGv{�h�F�s0�)�2�(�SM�����Ӯ��Y=ۤ:f���Z�$�_`sGA�^�ӘJx=�E{��	%��4��!B�D��'�dﭛs�l���Z}���>/�48��t�I.�*#� )��±b�%�*H���N�R����&�8s"�7�iEz!��B �~�o�T��̡�`�Ń�
���ssDSGs�H J�2�Z��3�<��z��K�������O� Fa��(Wr�e�4�JGC~��v�hH���S��?�9�(�Ͻ�-^�4A�k���E=찦ռ���f��:p@����~��۴����e������o H, ��ǏU��Dh�\g���C>Z��vc �*2�=u�3B'���"�� i�xL@)����X��
����b�U$�p�<�u��� ~%�T��3��+�c�1�M���>�Y�^Z�+�&笶r'֙B�-K��a����$��N:>����o�'��$���Ӭ��K�K��^$�#�|n8����
���2v`⬏�T6�7��ܴj���������>"u;��p�'.�שI�J#����*����5�]�n�7��͜����w(���cW�����w�O�	]�O
�����,��=��������˔��k��@�����ݮ����$��{�{o����+��Iǈ~N��&p����N+d�x�#��&��	�]n��ú�ETw����m�"����<EV��q�?ק�>S�g{.��M�!�%��:
,v[��v�9, ��YEMڧ�ԁ�rN�Y��/J@��y�|ؘ���CO�t���ޟg��?_v��z/l�zܭā1�㊮&�s���3-�k�����}���M�:�P�e�1IU��'x�5���­M�� *�̿�Nr�)Cs�%��V��arV	����N��XJ3��޾��*V͊+q4�y�X�3�u:��\
1�Ɗ͡?�f_I�2��d�ͮ�7��m�j/���NR�T [C�z�7�N�LXӌZ�4��j���2\��F��a�O�g����'���M] u���@��B�+�'vS������Wj��r��p#ꄍ�������`�����֐�!�@XY>��	�M��D���d��4�F�+ˌᨎ�T�gM��@�G��*��7/��n�������0��Ϡv*�$�L�Qzf�~:�é�HI����O�HV�~�6?QH���ݘ8������� �g�Q�It�%��:���9�����a�� �����Gj����ڃ�7��^�W�S�6���H ��(w����H�(9
;|��_��I�Mc�ƾZHY@�-o�%%��ɽ�g��o�#�_��y&P:��F��俨W0!�V#�u�� 7�)�������d�L$�"}����X��$�~u[��)���@GT��Af��W�s�Psǡ��A��o,6�T�"�β�Z�s�`Ha�er��TbH^�`$��/oYC��u����u��U�%<Ay6�13�]S�&���ު�^��Mm��� �NR@��(�Jw��!t�hJ�@��W�6�|�j���qa0W��߼@<��R�~H^��yQ݋0���3�i߬x�cB�N�����pg��,B���S;�5��!�*�q\���v����骊iV�̟�\g�H�r���Q�R�XO�a� �t��D)��!�;`)�pG�P曮����S��7��Ɩ�$�U]���MY ��t���M�E�|��J��<r3�����!��X�� �\CA*��Г���� ���
9X|L�V���Nx\C�*,�� ��(Ѥ����^t�����㿬��t�^�\��C��wO��Lf� ��Zv|3I��ƠRn�
3"�bv���c}d��t�u1 �9!l�9�?"�g4�O��^l�v�>�q�b
�'���*���^)��c���G��O�Y�u��������
:ǂѢ3��,�Y�⪹�뛫�%6Z�Ϊ�IM7��#l��#�s��S����T9׸]�4�7Q2p��OF����N�?�i,�[!j����91�P
]�2{����k:�1<&�l;�������fOU�||��m7�c�{� J��ݫ˧U�`}Ek[���&���?�s�����j�P��ոE�!WXIo�(	|�Q���<!���uSz���FJ+�N�CQr�u=��h��sH�w��5m�
��v�Y�-�J-� xW�GwGn���𴉄�n������Z�#Q��� p��D0ҭ%���A�ㄱ��B�e�5��{\(�.�'5}$�r6����?��e�8�|��_Ҁ��m�:���V�RaIʌ��^4��{��Nd�0�%CNǮ�a�9����UO���5,�y����>d$��y���$umJm3Q�ɠ�S6����h3�>����l��T����i�%��h�<�_���y��lP��^R3s�Y�Y���zh�BS���R�l`���U,7{X��Y?�v�mZ�I�[�70�E�;�fLP~ldHR
��A{���H.3�_W�݀f��I�{��N��	��v���
ʾ�h�`	���[���2�u~5)��3dq��U�ƺ����0Wa�"�U���$���s���HQ+R�s�ج��1�P25�7����)��@�],^��p �
"A]O3NPŒK@L��Z͏@`b�;��L��(=�������8�(��m/'/]����������|��Ӡj��ː+��qd��q�?�\�Zn�#VPF(W��$"�?A��+<ej	�%V�ǌ����l�ˊ���� �@���B�н �9�g7��݃l<(@.���"awF���L5#��-�h
_L�LZ-DθRMX���h]��s�H>y^G��=8z�ꓛ��^�5g)��w+k�Y��B:��=�lK a�����c��m��	"LG����`N��`�Ke�0�1A��q�����vv��0��{z'��_6Ǣ�kX��IM�.�͝0eS�9�	��%�p��
���ڄ���dE���mr	��19(���sF��V�X)�c��Y>���"�e��W��T�����ZBWTK1S��O .���3����y*�A0L��R���٩%�n�a'Op%���;�<��3޻S2������#��3&�jN�te��$HxuK�y�=ai�]��n,:m�/����[3�S�e�ڀ1;(>��}Cd����EN������q�3���ט����J�\�p4,m��@A��2�oy9�c�,%p�)��FߚTXJO|nw :Tw���X�^���	�w�����|� �a��#���·��غK�X3)}�,���J�yȡ�b6����d��J�*�=���q���0}�mAgˬ΢h�$�S����W�{Ra}{M�@.o��u�m��i#Y��Ҷ�w�?dN^X���QmQq��6�7\��<��*S[�� �����5�X��$����
6Ȼ�Uߚ\�@�H���mmS�{J#R��z��@�?(�=W�
�JH�=Tg��n�S�_��r��iAT��������m6t�=��K�>�f�m�}�ք��~�X�^tF�gq(�[���i�Yz�d5��r<b'�=�D9�x��Pe���nJ�D���D�Q5�/v?��Lo|�īl�Xؼ(��<���m��&���UΕ�Ȇ�� -�����O�23������)�~��rt��X��\��4���(� �G������D��Nn�#-YIZ������2w��z�[�enS���B$�nhh|��zg�qI��a�ce��_�nHU:�T2�"���;����ZC��5H5Y�IF���0Q��~�2�es���$>@�̤�$��F�ЦeKI�� �$"֪�����靾WCr���mZZߋQ���2o��h��Q�;�hD6��3$�]�9�Qe��ۘ��%�r�$�"�X9�I<+U}��{�q�v?+��+���a۽��z�����fH����^Nl�%�Q��$�������Zk������G�O�����B9y�=�.�9+�%z��emHb����ހ �[�IYJY�95	��N#8}l�'_<�۞=�����}x�EL���j�:$��(k���A�l!7�$��2�I�v	��fk��7��-�p*��Q�}d�5)��f�P.]���Z�����@���m�-F����[L�|�R��#X�\��s<=���@cC�������70�1�����(YNⰀv3X?3�N��u ]�ت)���8up]���Z�)|xѱr����,L�`����1��t��O��Z�\�N�DF�ˡ��?%�g��w�^%��0��6:$�λ(7��D�.ӊ��[�7�O.�����Ӷ���UO�A��$�wUU��	��!׎��s�3ݭ #����u��>ZYXds�u4�ziC8����p��Q>�M�q$����弿Qmph���{{���h�z6/뱷��#� 5$qR���I>��.-��
�(l�k� ]R��{kǓ&N�~����} ��@s���O��C� ����]�	���խl�3�����G�[h�?��r��>	��J��Zc΍J.Otмw��sJ��|�?�Ts����pX�����?�w����:#8���\m���#%�KÒ(�-��,����c��e�DWO��}��p�
&��ѢV��Z�([N;Oze�Ph�HipL���^�yw�>1N�����=M��~ª������x| ��ג�?ڿ�5/כ�X��h�p����!��i� ��a������@ 8�i���݋�h@����S�,�,��%iH�ٚ��!��m2	SF�Õ�(���r4��#�+�KG�����w�o�,��\��q��SfR�s�E{��6}��Yg�=����D�%?��j>KY��۠M�Q�J��`����m}�%���IXB���&_])���eg�1���V��jj���c`gi�����;�ؐ}tQ�B?��zy����W�2u	1�-�=��zb[���F=����+\��-:ݭ��JRV�"��K����a�v�I���F�% l�����8ǜ9W_�t��h��6��KwQ��h�{=R��3Ρ0�����C�!���Av������e).�L��k��f��7=�Q7�Q/|�zO����vud��AI_�!�d���M��@C]�r���QP�����K���I�������J�;�����*�>��D����-��f�H�7���b[W�1���ة��Ȯ�Wg�"��"k���Oxn�y
�
�U<;��p2�~)
54�Hz;����Ta�N�Y5�2��u]n��ָv|7ʣ��.o�U\�A�45eSK�C�N����n�&��A��c)E������������`ٶ8x�z���A#.bf��Kr+��02o��̯%��ln�cЅ8���Bp��l��dJ}�2�:�Z����AN����JIB���e/������*g�iI ��� ��q�����SK(V9C�4q�ql����Y1�h$��j@ݭ購D�$j���MN�Z��q�I��P^>Ǭ�-���B��o96��F]��D�t w�}�q�ǭ=a����]��=}^f��Bn)c��,_�n���ܗ����z�<����Lř疎"��IAiZZ��̿��(��W}V��xDAf�ٰ�[��%o�+M#�9T,���E���N��	�5`��Y  �ij����]P�U�;�[?��³�8p��{T�g�z{���Y�7̐p���ɽu�	.SC���{CR*��Q��J��S�7-�?,[���7 ��f�ڛ?������<6<�I�%f�����gN+�$���t����'�Vz��w�g[�E��ȡ��"z�0ް���+{;{�cV�Q�)�����gt؇�L�orw��j���?�Ǿ>��ΙdMr��a���c�e�l?U,��#,�U���f �����T�i���;pi���B2*�|��#)�{���#˛cp��a�f}`>0��?D��X%�ɭ���ÙIg��9�,/�hY�_�P�|k��X�e+���/� s�n�WJ�5ԟߨ����ꌍ����9ˏ�<��E����3.W�h�����0�3x�-$��g���-�Od�����,�D��:���4�����5�s�%��,`[��.u������S�+�klv�3̎M�a�и�����iKP��x2��GE�����5� K|���J��;nm*[�d��:dX$t���% �viPԇ�rܫw�.}�z�fsY����$7�ۄ�C��C�+��%�}�N�'�/НA��
ŹS3��>i��IR �*&%*1���7nF�ӕ9����/�f���lۡtp���'�Q_!g�ݐ}��=2�ݼ�*k�4�?ԷB��G�^���~�CcE?��n����ֿ),����V)�SɂCU�h��'%3�'��rV����#w	���!_v�M��G6R����L�.���8�hP_��lj,#���]n>�zCh3LNg�o�\R�;2��^�����@�6hq����K2S����Y%L"A����́��3ׁ��v��
����h/�gL6pDt	�\��F{/t�*KY��w����8�2�|��6�(�`���w/�V��A��5��?RZ�	�:�E\a��E�F
7	����G4���B����苕�ޥq�y�Fv�������{�<pF�~�gt`9�����r���f+K!N��H�D3'�Jm�u���[~b���#�L��c�1���t��`���O� Op�j)? ��vm����/��$�G���&����!끟�#@�e���0[c�k��U� �U� ���>B��I�y����%��z�"��cFFrS)��(?b�"����/��=�+JQ�ł�䆐�����J� ޫ��~X�t��L�G�ҬG�`������)�e��by潻��(��q�.�ܛ��9���9̑`�(;',�P���OW����+[�j��u/Z	�"1���ݠ��*C��P@��+&X��^,��1�E�fx�Nk�5S�aL�6���b�{��>��ab�p�i��nd̫���*cX霗i�c?;Z8�%��_�~S�@�p���� h����~��+�I���8ݾ�[BǱ����l�t;����)��pW��t�Q=E=Q/��^�����7�3=�'�g����mO��n�Tm��l4h���$]a����`T��T�%兪7��Ow�Pp�th��'��K\�!G}I=�t��zh�3�ig�_�^�^��̊hKZ����r����m�K�)��G��hҢ�l�kn�#sgl���o)����y��P����t�zد�݂W�5u���|�Q��@�/9H��NS�'.��'�Kզ�V��1�hp����)����H�g8Ez��t�����k����u���p���k�������k�b'V��3o�9�����l��_J�QS.:/گyˌ��L����<F�+0���VB�z��`6�.��|д�Fd����U��B,�òJ{_�u�/F"�<�5�{t��H�O˄Ё-��BJ�r5����V������5��@�v��m��$�[^�	E��N�$�����jv$�ů>Z"�KT�� 34.�Q�u�b�؛:O�q믷#�5�5�.�j���X���_}&���xJ����]�K�+�����-~��:�(e݁++�uK�cq��v���}���m$V���v��C@��Qm��NZ�m�'���%��K��bXƹ�M���;-���d&Bf����ԫ.����W�ǉYjo��|CT#�����C���v�,�+��2E�=I��E7��R��������5H���'�d��$�ҞtI��a�ơУx��y�LE�r��xH�ɋ9�L�ە��'@KT�p"���Y�睱�t�~�����g5���N���?#��ܕs'�6U�!��[��Ӧ.�"(�t!�������I ���#��o�"�C}p{�%�6�����<kQ��u��ɠ�������EV/����~7����;�k	���Jw4i��ɴϗ�H�	g�|ٚ����H���m=s��M�
�ar<scGs��]ד# ��N���UQ�)�n싫�;�z�e���vH�P\�&���"��R��W1��q���i<�[U�����<_����ɔt�sD�}�o&\)A��R�I�:��~��W^ݶ��
z���p�=.�ˮ�Ʉ>8��5V5=���K�9J%���2͢[�k* HO�&G��X�,�� ���;���T�@�~����@u�S��~`�W[��������Q�vȁ}E�_Wr �������#��R��,���(�GN����R9���sf��GŪ��Ϋ�H<�f-�%w��no.�bܐ����2ii�mp=�(�3��f~�f����*���v!��ldHw�G*���%��`��x��"�I�Ů>-ؕ�R�ɘ�{�����d�	���l�˂?�u�ӹ��5�R^��e�O3vb�R-����҅�hj�\�,5��� �N�����i��ˠd�O��*�lp|Y�5����1��cc`..,�l(>7����8ݥ�q��rD�@�.�[��뺬Lw�OMs2�Cp��UTa:����8=?���L�|	PTWU�,�4���` ����:(�;�������:tP��������^w;�_�Q]�	���ֆxN�zs@(�8h������ y)T�f�ը�M�S�AX罳i��h�jdP��EЭO�����xW��Zw0Y�ج]���S=�����!6�3I�Ea������g���s�
�O�M�B��� B��?Q�V�����K��+c���%�4x�:v$�с�$�Ū���c��V���=-�҉G T�E��"��� ��$߀t���b��efZ�'w1���3l�I[! /�2�l�a>���a���1��N�p���a���c:��c�T[��u�M�d<PL���6�!z�HP��й��E��#���#D���%�0��9�SOϛ�{��Ӫ;��	�d�zd|�ϊZ�|�93`�9��%�����Nƞ_-�slv	����O⫰�_NYh�E��������G�4�{�ld9��Kc�%1&�v�n1f ��#�m9�d�H��o�?�P�?R
L�Jӂ:�q$���m�1Ӧ�p�pS���Ą���t"�c
ۀGme�Z~4�o��h�/g{�ƽ�lJm_�ˈȏ�ϋ��:ÑE����?r����_��WE3R���N��w��՗��T6úl���[=�T2:�m>-���M��·ى���a3�H{#b���3�K�'���s�8[X���6�M��e���S�	*u��ϓ�s|�L�(W��u�a��OA`0i�Ԝ�����۔A�����3H�� ��60�%��z����y��������`���y���������Ѡhax�P�8��2}te��Rˏ_�G��#�zC$(�� P|:h�QG�Y�Ľ���~��w;��`�|�,Vx�"�Z|q: �����r͉H#��ղ�ƶ?\�s@C^!Ǯ�."�V/G;$�	}��
K���P�9��Ʊ�rV�]��3����~��y�n��>΁"K���(u��'���,��޸3�F	���6���}{��
jq@�)P��A|V��zaf:����;�c�$|c��� ,�k�޵�&Ħ�������*GT�~hdlOi��5Ǻ�� X^j@�K�%���e���T=x����}HO�XܝFuJ���8��	�`�w��`��0��g@�m�,u�*W���f�������-��Y��+�S����2�'Z���jk	��"<�+	+Wwƽ4�Sѻs���a�*��9b���#S�U�)>|�f?Zp�'Ե!O���k��:Q��{	��hT�l��aP;�pB	��*�j%���Iz�M�J[��F�nR��C(�����7���]z��$��xP���	ݯ�$Ll�� v����y^��E�Qg?�V\��AJ'hW��ۥ�u)�3����sJ�sǇ�&pm!������Y�Ɓ���T������m��Y�ԃRD�ʡ���4~ӿD�Um�~����*@H� �xcp�⎽��9
���J���u�븄svJ�.�vs������s��O�\�h��%���BK��țU߱z�IYd� "ς��_Y��iE�˓�c?�����^��ʸH~���V�-A�����r��Tr�n���z;�<�b�zo ��*�	s���ւK��h2H���а)���%\��/�u��3��Z�������J�m�d*��v��*��qŰ�Rm�>�O}@�Cyb�&��֣��=6,\a��͈�/�C
��
ù��:6�|���B�Q`��{�~ߜ��ځ�f�n¯�s�y�V��wqko�
*,TYSלK�~���1U�ѡ�=�����9�I�ke��?��{�O�r2��`�%m�S�u�r�P���������(K�iM�"�o� $s�7��[7����Ů��Lq<Y��K�ۖލ.T3
��ͳ�N{���./�ۧ���}l�7]-�_3��%7»7�i�����j�ӋR�?H<�1��.�(W+�2=���1A�xh`���l3/��ő�46\���tR$�+�ߑ���Ma{\ɥ,P�N6i&��
K7�T�46�MB��=�6Չ��$T�Fߕ���GT���J���ر�^+�)��CJh.����j�#�pT�B�gʇg�0`3��^��K.��M���x��P9�CNP�p�-x0�����Z�S0>@w��%m5#^��h;�N����AԎֆn���9r,��7#�RzD���U�:�I�{�����rz̄=�����;��� �GNB�mm=��7�Ӄj�m�ߝ�z�����,�}�_��/�*lq���L�}���*�^��+w��wG�
$8��߳� ��D,��<�퀶���{���	��n�����t���N����w�Z�T�W(A�K�*��#Y��}d��b���ޅP��Y<ԕN��)����l�ÿ�=��Mu�{R���IE���) 㷴G�jc��$�}+�_��IFg;��<��6.��t��gG�h6�h�Jc�$���_[�D�n������J�W�%{�7QQ-]�}:6�� HN��E�������������<͓�f�o��q�~�:_�H����!"��齖y�_�i�ŽTL�����ڱm4�Nf�c�-x���k��0���lN�ȁ�-���L����.�$˖��L���nB\��6	�W+F��܊�g�G�����'2��=Q��W$FH�u'��(I��N~�J��8U�\�0��$el�v"��Ί5ѤT�4S,�#!��d��T�����a��k�Du��P�mg�JD��h�@�ڄ����
��	�>�Q6*;�S��;H�|!-VE�d�S�B��՘�&��4��b$[��̵����fJ&9��C�.p�x$�5Aث��"����5b׍�*�K�+
��Qy�s'���πw]��S��nC�+5Dդ����E�T���c�5�6��1�`�|wE/Kȇ�g��_�d-�a�&2�e)[�#~J�^��z�n���&TC��S��dם�D����(�w���\��t�?)>9����n�iם���o�2?i��� ��Z����Cw�e�΀C��}��.c>����^�|�c���o�R��'l��v�6
:
�&���\��hf �Zh��J�/�)ܦDBR	;��'��=\��,����hQm�x��E���c��H�.�p.�+�\�`jj��T�m���@q���i��2J�F���d�kq�C�wsNġ �xc��S�Vv��Y�.>D�C��lX�6~�Nu!���4gi�v�^���ru!�;�nZ�bаg6νH�Z%$��̣���Bd&�O����葬Y5�*�ؽ:���b��ˈ�jh�
n*��"���Vs���',����3�⨈Lx��4���j�:�Fȡw`�J�d��Exr�7�vy�H�Ƙ����6;p4�]�߲`����ۚ� I8�Y���s�M�c��n�@Qga�=S*���ݖt'0Ӟ��m�aT�9@x$��Ӻ�3�)4?C%��Q�(��T�S1h����S��P����;u�{D�<�9e��rXK��0�$�t8�:�9�A���<}���4ֆ�j��h7�ha�:�D}^����Co�^��7�����|U��+�'�
�P��a:���$\^_b�=�䕰LyZ(�&�ԭK<��8(�&>�n��uTT�e=���5�n�4ϳ#4�jv��j�H�p�"w|�~��	�������`�4���#@��Y{;���;�Z����v��s,� ���ρ� �����6υ-`2����7Y��x��%tlk��m��B0��SC��c���v���������=:THE=K߂����;k�Y�n'��D<O|���A7�O�$��Z�����dsR�7��NcF��ni�6��&_���{m�V��*y�ǁ VNz[cp�v�$�n1�4�uT�N�8����*�|3*H����1!
��!@e���������e��T���l�Q�Ei��?2��.\ݦ)����	��_�|��� ���b���d:J��X-���y@S�
x
k�m."/����/�ވqع�t��Gg�IB�[B�C�jb<����U#ǵi��a)?�݊y��\�f�5��>���R�~��М�Q5`�3�oк���(Q��,�-�ћ�v���%D
�[2�J�ѭ�+�3�wۗp4��|8�}���#�k�f���$��U��:|t�t[��i9��~Mɣ`#��)`��M��2��ˤBD�Y4>��	�D䝣cg���}�O���J��{)�<�3����\��U�јY0X�&���<[/յ�Re�ޝ��Q����$=�vBK,5Đw^��Ƀ4c� ��I�E�BwT�}�V�Y��{�y�� ���'`��������3�6h\(5�t����6YL��y
�
��w,�7�-+H����O�)�E�����K�[�dg�Qo *�l�d>�~j)b�q��71��#]��8Z�
��־{֓�u��t�MiE���OЫ���3��S��'��ͧ��G=�I�rl�%WhS4@F� k��W߅��N}C �BZT���~��� ��z|��^e,��v �}׋��`@�&޽�r6�8k��v�6@�nS]K��z���X�hE�5�lK�̠$|G=��9O��^��N� ό.gU#�RN>âY}GT��3�?�����F����pU^�pq���{"�p��b�f�3v�sK�}�T����_:�
Kj�'��m�Zߺ�B�%��i�ִ��'��w]!��.x?���$i�b��z�M�#_�_���Ϟ��a�̑��� %'�C�/Rw6EY�u
1�K]��n�f��G�H���3V�G)V���ytH�,�Ҙ��t	֖����]hǱ��Aa�e��Aőn����"��)���� E�iL�#���I�����ˑ��t�U��g~���1����­�$)\H/����OzS(�/�8�����ɂ��wi�O���G�D_h@t)���*�0� b�xXN�"ғBuB���Wp��]Z0�HDM%�y��SX8�v�� �����'�� �O"��c��,�y̬�����-{%��9��� �o��-��)���:owd��E{7{%�9���|��c���x� w���p�2�(BB�W�l�E��Dj"��y��|�k_���9��0��U��_�h��'5���U �e���5��U]���)�>��J�P-e	��aB�1��Y5�l4��l�š]?���fU]�<{��E�(�����K8ǀ>�뵡 %@�Yn�����!
�KsW��c|�%�"���Q����hz8R��x���y��uK!\��*k��O�%#O�q���M�����d��O%�p�z&����ޱ�Q5o/�W��4<9�U�~�-<����"��/5N�b�I�tX�m}ɡ>��e]�ٓU�=i\�P��J� �p[C��L�v��\��/�YW�-���s�5J��z�9��(��uWГ8�ti�@���e�3�J��GZ%n��C�@���!C!�M%�ݻ��kn���n����ۖ����x�d�x�UVͪ���e ����V!����}��	Ϛ�瞜hUi��Sn�?�����]��4��n���է�[;�P��G �K���T�p�O�t #.��<�V<9 �I>�P����"]���R�V��Y��z��R��0>��1�=2�⒧:CA!M��@C��}^��bF@���MY㝂C�`&��I�lU�#>����)S��ms�O!�~$�,������X��a���՞��� y�%���M����ۍ3F�[΍���Z_���B.&F��d*�놤��Wȑ�@u���틄e�æ���+���D���W�c]�[�B���y�wS���/���̕���U�]x,UCp��;���}��s?������x��8��'e�8"}���Cm;;`}il�?��cnopm�/��!�el"<��܌���W���f��n6��S>���&�Goe��_�A���'k�����q�~����C(0�0H��
�E���5>i�	N_#Y����uɿf�"{l$KOF%;���<���'J7��ڧ��ᬧ�t(�qe�(ֈ��c�i�ܱ��Y�a`y�HU�rǣbRt����>�wo怠�hC��7R�-�@��Lm�LD��ո}w���☼*bn*R["��*�� ,	EF��f����r;��z"I��BI	R�j�ZîX#y(�}/�7�*�Yt1�Q���	L.�\=��D;�����6(�`~ϝ9
���=�M�ZZR�0D�7Z��~�ff��+@��Xml�uCAZ��
�LǷ�Y��j��

�G��9��J2I-�?�i�����0^�@���:*�����i�_�y�!G�y��EKN!O�z�zl>�����|"�
f� $�gn��/�����x�)��9�`��J�ak����{�����;�/(�߀G^D�k�Cma��uK�>�/{�4/�N�x�Ul��yl��u������J��4U��t����?��(=�'�����I���M�Ы��&��Z��:��?�V��n�!<��֭�%>�S,hR@#�����r������.̂HI},L�8���I&�hhN�t�j��)�{��6�`ζ���Y��<suݽ�~�p��幔�������	��)���N6�(`	x�x�l����Ƴ[gl�Z)Y��EF�7 ��,{������O���9��k3o��@�/o�Ve;���p�k�8k�20V�&w��~F��gL��Uݘ��,�@1<���ϻ�RjيMmx�jY��*|��0��дj�e���/_�E�k#����:/�ۧM����$`���(m�f3J�b�(��h��d�Y"�ل�-vANY�T.�]�&��F��K�5v�m�(h�w�Ť����5�+��\�D�����\
s��^�8{�,��B��Χ�v���K<#L�=��#1�o>�`�������M�����!�ͭW��k�3�D!��6���k[��ɜͨ�O�s^B���XC�i��~[|W�Q?�2k�ɹ�� ���@P���m��-��kN�w(7�f��D`��� Z�>��cw�������Oo�E�p(�9|�ǲ�^?��O=� �E��Q�uE����� \2�;]�1)��u����`��:�W�W�D�B8�VX+�b���"�Z��Ȍ����Z�����[@�|Tb`b�	~� ���}�楢�G��
��G��_��Y�.�.�P�_���@��q���at�Q�F�NPtջ�D��  [�2�S4a���w�Q�]��N���NL�in�lw�2�>3��K�~is�-c'R:�U�5�/]ʅ��Hrn�zS1F.su}����CzW���Ѷt���a�>�D�#���4$�c�4�d[Uw3_}�Y��m�	^q�����8Ch�O��ik�w�(%�-ڌ�x���S��T����"�'X��l�b�B	�Kd���_;�;�I��Z�kN.��K:˄���Cn�nW���>e����������_l,���P�׊~���+ Ы3������W���hEnZ���"�I�z���{��M��W���~��Z��U��밢����l[L��q}ܿ�8��q�Ƃ�M���{jaht.l)��E?�������a��lc.�9k\�dp�&[�v۲��R��qA������G�4�>�"�M���J{���b*�U����?��� |�7���;�)Y���y��9m��Wk���Ձ��b�<��~/xt�q5����2+WZ��X�T�T�벲��lBF� ��?�l��^=�n6hr[�>����4��2������j�T�wI^�ܾƌ��jd_j1��6���Q�U��*�͑�6�Ս.�b{;��B��f�v��ņb��A��n0��M�܇>�3��OR!岻�8�(��߮��"��Cj�_c�b����TR���yx,f�U�s^��i{κ�8Gt�x���U�_u��� .�I>th���	���FnxT��1{�ސ��Qāt.����6�U�>H�g�<kO���i�{e�F�*�A���;���Y��p�Ru��Y�ABC������V%��!q� �D���L���Ge"�����h-ir�1f ���������4T �'L�o�i;�����G&�\�r��Z��@���z�:�� $�~�#љ��G*	�zn��bJ�9�+$̀�^�2P�]�-GyD�P��t���_[?kcד���qi519�Ό��*�oFۊ��w_� t��f���:ׇ1��:g��f/�Gvxi��E�ZPGqV�j��ڡw��}g!7���{�<g�Mp˙�<�K8ܨ7Ծrp�o &6$���@��d �1�%�X�_�}/>�Rl�
Ҫ��&���)j��?��L���O��H�X%E̷�n�w{q�!t16|���GiQl,��\�[my�8��#�e<�d�r��?ظ|̜���l��Y��3#X)��g����~w���q�/Jn�e>D����+$h�sXl�K\���}��p}dwh�iԽ�o�4c����Yj�T�Gݜ��@E�
��sEC+��x���MN���ؐLa�<���<�,������&Y���� ��_�@�Z�"kVa�RvL��G@ �����gGI/�i�{�Ov4�"�,��ƿ�菀�h�P�}j�32t��B#��ִi�e���v�P�UgT른��ZMM�(��ſ}����ۈ�qܖ�~��)��XɫX�}!'y��7�@��T�u�w���Z�T��o=�@BX[��z��Ȏ��]�-��qIK�Lۙ"d���uR��3�v��+:����b���*�M���ŵ;�sz���(ٌfgu�D���ds�;���V�KK"�@C�O}ŗ���&ڽ��j�3U�C\���]�En��J*��|��}��j��+���/8�2�Dmv��U���4�;�!ض�<CF�3��BF�&f��] ��L���x���?<$�|2UCGpC�{��i�v�c
���ȵ����vf�!s{4�I�K_91��P()���I��o�3K�K�{�k`��A<bZ�R���M�%�@����U���_��OȊ�,�������+�~^��� :���.�S��9�.���L"�-L��ɷ�s��JU<�����猕G��u�غW�=xL{)��h��R<^���1:�H�0�$��K�2�4�IΕ�"��M��#b�7~�5��_@����i�&�zb`q͵@?u/��C󠢍׵��+_Z����O4�P��X��`�6@��CIM)e0��둩V����$��D�3*y`⺚��;�"Aܷ���/\)Zn^�ܠ�8�����	��w��w[~܉
�_��X���o]��dGK��O-���4�7�
.`�t�����h�s��S�h���uA�K1�Q�)��0c��i��F�B�1��;�<S?�'��s�z�="�k X5�߂�P�n��T|H��'q �k���B�A�ᖹ����~Ꟗ����፿
z���O�d�u���#�����Ă_�W�5eF�4*�`-�̀-��jb6@���+�/�9�g��!�V�ۚ	�S���Ԣ���}%C�K��(�܇�rWy�`�4� �M���f�l�9��Ps�!�;-x�����,�}Y�:�r7ա`�ٍ��Ʀ�j�NOp�����& �m��_���S�Z�
���o����)�֫�I	�fL1퓇�5_��ջ��H�N{y������7�/N׍�����M�vm�q�!q8&� ݺc���)/~�g��@nϰ����uR-/Y�dY��d���q�ў�~���UL��-�j��k�T���
�e���x>:�hF!��{�úڵX��`�D����$E�?��#���q)��w1Y�{L�]�m�壱�^*S� �U9���v��G~S�0�٣�){G�H?�N ��6�4�̱7��!�n�g��Z�7�\'#R0KK����,���'��ބq�,
�S7�y��]���/���dn����>�鏅�e�j�)ՅzT�Y�)�l]Ѥi��M��5]+��QHF���Oz@nn�c$d���'k_�&���"�v�iK��i���!V�J9�2[�2O�+D��+�%ꭾۢ��_�M��u�-������(:�L����旍l Q����z��O_�^�4
���ufz"�cQ��Z��t�74KD��).�
p�`-pqv��'z.E\n�� �=�q)�5$y����zL(���Iۢ�����i��ڂX�r7��e.`Tğ�[R6IW�nN+��B-Y{���CK��e��F���Fe4&$MW�[����_|����R�/!��b���a���D
)w(�Y�V��͇9���0St����6Q١c\�6	�`��.hQ��;D��q?m��~t ��O߬�*Ha���>�S��<6;�Ɏ���J\�l�����u?�#M�$��8�lHv�lo���T�uj`9=_C+%��C����7w���ۅ{��w�#֥l�¿���e?���oEN��rl9����w!N�Ɛ5]_l�c?%�w�t{&����0Ee�7��z�A����S���$���f���rT%��� 1��z�C�9n�`�kL ^��0�Mj�.B_
D#��Q_{�ʮ$;h�-_ K�wc�	c&fw�uӬ��7��ۖW�L8��_W����.K��yA�U�Ǒ�D�1��yO�+��W0�>LD���LlWƊw!�<#)/�6��D~`mLz�������^<�����$�:6���%�Hg�x����0$�W��G��&7r�qRq������H�!�.��C.��)�@���`&����&N�����͇�u:f�+����V-��dT^ITU�z+�Q���h���߇�uF<lꦴ�$x�� ��=.l^����v
�-�X�S}�;�ȗ��8W恹�8�S��<W���Ub�x����h�A�em=ɦ��D��؏2Yb9)!Σ&�g>�v#�J��h �I<^�/�8����ZAhhԃ�ds�Qy�v�E:�%[�*<�-�o0�y�yBQ����J������jm�����q�1�w��/G){����,X�Oe{�'�/h�L�٧�/�9�-���y�Z�}��;�p(����v�×��cM�p1-ˉ�_�Ca� ��r���|�Q�8����'�,쭒s�����;�~!������h��X��<Ω��Wnq�ϗ�Q�u+o뮆�ce}=�w��)iJ��n�DxQ�}��ӡ,���(�G2v*s���Ѭ�k���,78�ax6ϽH����@�IJ8�]�q(T�<ԭT���e��Eݝ�\w#�9�
]lY���B~�Chy���ɔ0艬�X�F�����G? 0{3�YU�>��>1�1V��v��əU5-~;�U�U)�[ �>�W0�@֔�HÔ�n[�y!Ү�^*�&��B���� �pΟDn��f�����tC�"�r���i��t��I*-��ڑm��ڭ��m�2A �γh�Kq�����t�n*:�s���
nF.�v�ף�bU3��ubWan�*J�qZ?�}g	�=��y���Ȏ��&6R��DJ����/�ЏyXL�1 Z2��y�h]�o����4J�>�jM�'���O�6���)��8n�� �D'��@���m�MO��.f���'3����(�&K��G��'o%t�XU�=��1lw��Q~��[m�=���H3Z  7ߴ��h <���UFk����Z�? Y��h�*��B�X�F��i�����֫�OOCת�8��
`���k�[7V[FP�&��?3�e�ͥ(�O"x��2��[g���6CzB�����I��?@�M�/'��%�4��� 3X�p�xO`=:�d�q(%��]7u~�v ��^ �����NM��k�&"d@��*U:hlD������!�̵y��չ�6�6��`à���-��+[����l*F�[������S�c�W�1��M��d�x�����vaq_���g�4
�ʃ�j`�{I�c$�3�jċ�����Q�.ު
��8��{h������Y���o"�������b@�S���!�i��0uπ�'���P�[8hIUB�I��X�� �^��}�~J�5�����Y�M���&��!"\��e�{	p���b�ip�L�О�/���J�d<21���|CS��W�<So|R��C2�j˔���}+TV$3���x�!<���� Utxe�8ܵ��ĝ���_�0������T���`�T*��z9�U���#Q�Е���Oj*��>��*V�FX����m9�5��S��"/���\I��Ld~�}�xT��I���H۞Z����̮��b��DjC����w@fK%1���{Mp(f���Z�"�C�3��TFK���c����:���*F;4u@-���|�� ȸ8��B�m�Q�� ɡ��r{HǏ�8��A�@&�}@%M�	�Қc�Ȝ�H��^M��<#��]ȼ�A�{�>����ع��&c�X�����v�����L�է{��������9��;������"B�#
Q�I[�2�$.���I�S��Vd��}Dc�{�Iu�0(є��S����_Hڲ?*^�q�7��;�>�v���2
�Kv\Ɋ�������wC���'+���Z��I����m�hì��S$~���Ɔ�����A�v��1ߖ&��Vy�d�=��_�2&έ1�`�l]�z��M5����6��~;�#�Pke�T��lNw�/)�7�����x�6���Z�b��飽8��w��aA��Dr"�E;���X�B�uC�׌Eī�̑g�o����H:�R�\7y�3��%}[�B�h���?�1�l9�Ecg����^�p7��V�g�9�OD�t�,�+����Wj����wʝ�F0��U��uܥ�ͷ̂����`��*����1Yu)�흹����� ���n�ln�xYNj(�V4�]��:-�^�ڝ�eC����ހ�����I��Q�rm	��q���C�6�E�����f���Cv	R>z�a��b?�(ԝ++��E{�G�l�`A�*k�5��8<0��$H�׬�\|��v5���Z�o.�����EڃcRH�|��K����EՖ4���ɡ1ń����s�,��,S&A`�!��^�u6��z��o66�X���E�����T�O�}z�v,iE����.Xi�;fbY�
\��d���h�EXCz�)/w�Ђd�ݍ>ê�a
��A�d&frj	 ��)"=0u�Ӭ����o7�\Q�EB����;"���F�d� �m��)�X�<��,����#�v-v�UB��4"-\�r<�*��Mfϼ�;��9[�C��.�Z�Ro��V��e�3�(��t�k��D�|̋YWR���ʄ/~�Pz���7t��F��lT��]�'��,���kA�U�N#SG��P6�ĴV�P&���B�C�ڽ��R0�K�vڢ���� ��&Od���i)H�e^3Ć��WJ��JOJ�4�����*9N�Z�&p�76ϫwBp>�]�6��*c�Ŵ{��1��K����ѕ�M���8S����Y�N"�?�X�͙-z�P���W`'�I�����2/s�����0�c�������XZ������u�A��wzA�g�$b3}�m97�U�q�������n�,I��Iϱ22��V� ��*��"��ɻ0���I�	�ka�y��	���g�$���SVX �Z�	�:����;�₏�(P��`w.�����n�J'���k-UKU�����bI6p�10��"������K��o<�b]&�0�i���3�� �'`�΍��MK�^�==�1�Ik.��|�I��2�ƥ���)�v�d�*�S�a	f..��1Q��d�v(�nr��.bd���(��u� �v6�d]7a���sx0������36�����*%��dP���A���_]�o�J�j�f:=N̜��9�|.j��������wSKA7a��O����&����;z�ِC�vڌ�'9N��	?/��W4=�s�&D;݁��L�[�P�J{�QR�j�`��6l
3sm�f�����3�l6�E�����Zl��mH��U��༦�oX/a+u�g�	bU��U�
#����"���o�O�fj��&=[7�8P?�ڇAR��mG�FӍz�䍋�T��2�91)���'�qoI��]�{W�GÀG+)��Sr\�0N�pgOLJ�x��D"�Û�bۨf�Ƙ94�̑�	�π <�S��&E���9��L��,��US��2T����e�/YTS#Lwd8����W�B��ύ���fF��K_�
yϒ$B�"��l.%C jJOJ=���7s��j�ʪ};��ڪ5�ޔ�Z��Y��[
Ӆ�/F-eC���#��|KrxA��DF4Q
Q�E�����ϡ"xI��F�μ	��_�Q���s�Р��G�i� 0�9��:eE�t;r�*��t�}���i�sr�N ;�Aq��pj7(�E���Mc�c'�h�a��y��u��:eg2�y ��-2>	%HYn���0�|��N��G�����B�-��h5�������h팱�`�/�ԓ�߳�qN��{�x4g�������Vո\)Jł���Ib�3ċ��d�\ikM~Q�%��A��ը��@�sm����PQ釦�ɢws�x��]���-�Q26s�ap����-3����/�*�5τ܍����?��wk��;蓫6G�_���R�}��T�����O�?�ep]��σ��ݽu�m�m�X5-0�~ۣ-U�@��1t��7X�X -��x��w��K��,-�7O!�W+Qv�"l3���gAU�I�dB��o�C�^,M!����e�x�*O��7�x̐�MM('�~`��D�l����.�i��p��N>�}�7���=�l���W'P\�K��v�#�"Nl=L��YA؟�ܔ��y}�����!�K�Uى�$L����
�,L�*;�)G��K')Z`�7lW�%�׿�+��G]���3��E>yŬ����j�EN?d��
��r
{A�to
�ro���̫W.ж��{�����S7�<{��w�QXL����Aꁎy����݉I~֘���B�n�&9�x&�ߥ�P(A�d��;٘	"�g1��������t��zw�OL�.���*i ��%X�-�r���Ep9������R|��?JT��������|>�u��������;����+7�2��ˈ�D˃�DW��71�K��xCn�E�+�A�D�~l���R�;x9�9V��1	�Dc����%���|����l�"�:��W�mU���x�����H��ٲ�Ҹ��D�~�K��g%���{Z"���b�X=����0C=`:x�z)�h���=&OW@�G��b+hp �=	�c�/���}�Yc�1�x}��C�A 
�#Cȭ���<�]�L����E+�wa��
�3�;�w��$�d��04���$���˹�=�����*�p��|2���u�z�(��@�L�7x�����0D]d}nS#6n�o\Ù�u�Ԁ=����b얢��좸���ڱ���v�:�A1������"�ǱVg�9R|�������f1�V���劈M��^6�����?r�Z[�� �J��y-X<qD��ؕլ̻��W�2��<��ԝ��Y���s�E��P�8��T�*7�����Z��~ُ�"Grg��e5�����y�k����Y���jYP;A�g��o�A����?T�'��fF�"��N+�����U�����:&��8��FB[����Ua�_J�ܸ�N��)���EpM��I}��D܌��4�����O�A;��U��M�Ӛ�6�FK7kG�9+��Q�����NMb�>'�"a�qXy��
6Mܒ.ub@�/�� W��[	���ޕvw�<tc� �"�F�-L�b�Իt�����˛�N��.��I'y^[��i�V��V�&�Y	CK��n�������Q��&_��]��&'�U*L<��M�J�l�2��k�^t�;05�s���l|�E���%�5��-X��\@;߹�Q��\%��)V��VV�yQ�X�������'^�wh�������4M*0e_��:��=�
�I�.�We��r���'���"�%���A��"8.Q��ÉX�1�o��u�(�1�pzQR�+5��:��D;O�f�I6��RA��ة�-�dMgȃ>�|(GVu'm�Пg�fgfэ)�D"X��9B+y}����$5�Ne7Rp,�:�C8\�<�^�u�_�|v��io�n�R��&O��o��dyޠ�Y���-,F�&�@�-�,�ا�7�X[�>%������*J��܁������!��S$�yCh�<�y��O�{��-y��.�*��;٠�P�M&VB\:ҫ��p�uȦ�>5� ;��FT����v��0Ӕ�XꨵN�^-���s4'$a�2]���gҏq�7�u�6둳R��ʘN����� ����nGp#�h'��%ׄXpn@]�c<���*�=�`�����ۆ�Kn��T�R�"��3��WDZ���MC��C�t�x�|��J
����V�M6��;�95]�a"�ܣ&J�f-�+[�=ՙ�GjUK����I�>�&��x�Kce��P]����l&c@"�X�J�4d(�Ac�FNy�D��4�ػ�
&e[T_u�k�;ɎFZ���hR�O��8�#�$1���*$2oِ�� ��(�hcP�@Ե[I�;���V�P��'�)I�}�� ���$�
�X�n�t}����i�>F./gWx8%h7�V�5j��Q�73��H]x�
�O~�f����(e�նOL3��DB�6<����O�a6� �(�b����`�M��(L�񲖛g��T�)�o1Թ�&���d^C1h�#sY�
����Vm���Vv#l{�i��G����:O)Ǝ�s�Y3%:��X`�UFk}&d#���g������գ䗘���c����@�a^���h��YbƠ*V`�y���� 7��}��Mn�`�ul�1<���-L�F��[�$Ö�H1�8Q�'�o\�/��y�4;�k�{@)]�/�Q��|Sc��U\cN��VS�~�v?;���nT�c�F�?���|T�x[�|=�Y���5���~n$��*���Q�*@�#�!�=|g�&�e�oG�� 7��
��h!C��Lo_��SX�9ΣW#���g��V�f���F0��	s���N
��ئ@�iQ��0^���n�JL�q�uv��|�Q�Y��lo��ojH]��e?��z��`�����`�#u��n#�O8 g9�oo{�#ɦ9N|�on�Ty,c�A�R�>���������fؐ�v��7���`B!�����2ɻ���Y� ~�ru<�|�{Y�TV[[�<���b�?�p�T~SX�cBn�&�ϴ)v������U-�X��D- �ޘ� #��<��"w��d��ki�hͳ$蓍�H�w
�̝߶1mfL6�*��qi��,�u�!��vTYz2���
&YĞ>���\�с�C��g���9#ԃ�>s��J^�6���ͫ4h�e�*vn�w��{�0"Aw���;AWF�.�#O�P���c-����!k�������׏�U��d��[Z0ib)5�{�=��Y��<�LT���l��f��Y����W�B��UL3w�Ҕ_i�7��j	���舡��3�
p��R��a8�&��� F+�8���$Б��J۞�E�D����z�C��v�N1�L#x�X��5oT�%��s�����5��cL:l�� �S����+�+�G��$�T/[5!�NʔK����H����5�ڈ��Z���l$&L��ͧ��#`���r:>�?��2 ��� U̵��s�#�~I߯/�^d�B���fv�6�p�L��l4-����
�8��\�dk�\u�̓6��Қ������������R�L��%�V"B�G�m��;��%ډ��?�k3}��C3�G/ɸ+I��^�5{��w�u�Q��e��Owg??��P����P�I���X��s�\d���#1�"����^q��C�A1g=1GI�M���xA�&���*� ���"A�4 Vb"7�`�Ap�w�	}��wOя�Bso!:ϖ/;�����hα���\��ￌ�[S����� �����$]�k�?���0�D����6�Ar�5�"�SИ$�(?��\0�������~{��� ~wK�����r[C"nNIа/�����~w�a��~�����R�
��I%</�5�G�D�<8�n��G�V/�� 4��L%�w����ى�:�o�K\ܓ҆��ب(�2�g2�&}U��	֡o��[�J�T(E�@0�g���i����8(	_"4|���+�%�&��㔖c 23��޺�qv}_�?��ڄP7��Y�K�ɨU4�0�L����>��N�UK������N�x_��)�T��D�����-�值���)���/��%�6�Χ���:e�L���0#�V�[�x���{**RW��U+k^x<�[f��7�l�}H�g���CZ�>��2L��p����9�唵� �~M����}]�ܭ�fM��Y�a���F�U�E�YP�Y��M��&�o���̌��a\A|s[c���:�Y��<�] �lpZ/m�W{	;@��4��*���W�0YϠ�f��U=�>8>-�GZ([�#� Ͻs'[�{
��M����Ԡ8�`��́��.�?|�~\@f���Ğ����*��M�X?�����7y�ћ@�zIR-����~ks��e�b�@ȭl.b��@K -��n�+�G3o5K��i�ڈ�G��̦%R>����E�I����l�4�v��B�������U����B+s�{&g�f����t6=׹A\��t�������r�e}���@����f�%�Tu�sOX��kƉI)]�8"%�]Wl�K�'y,�k��g�.ze�:W	7f���ŠY6����Ri^d����;�[N�:R�5b��O�c��"����G��5�A�6��y�+����:=�v�N�.��A���:CV�^|�B�r ��џ�}�)#�aqe&u�=5��!k�65�/@�^_�&6�wxϱKɦ��|�$N����|[[c�Ѽ��8I��2�c�_$������Ec�m2����K�yA�=�+b�nS~;�������F+P���2B�D6	�07�jL�6/z�8�����v��N4
:]���TRJ��;�K�01�:9MQ����R�*W@f�"�.ހ�xȇ���7������?G��_m���=���5��z��S��<SZ�hM�
�b�����&V'�vh{�^8<q���VR����%DR(���ݭe�a3M�����m�N������瘂�b1m-t����޲4�b���킄s�o�Gy��}���]������7:�W�(AS�O�L�W ���;ń�h�ۛ=�������k���J�����g���m+��׋�6 ci�ch�	)'�L �S[RҠ��W(fč	pMmRW��`��p3X����ۏr�ʭ3�J��Cì+@������v�K�LRy6c�("D�w��A>�� ���d������ylI����n��\*7�A\��TJf7,e�տ��}�2�t��7��~��9������POʾk�dU9w��DҐ��x�\���vb}������$Nw�;R�i�l�z�Ǿ�w�D��)_�X��>��8��A6��61�K'�(d�(�*�j�^V
�a�F|��ɉ��("mA�m�ؠ[�BB�D���k�:�E�kFA��M��	m_�{<y�p��7��["�����t����a1�Է0Y��AW&���c���Kv�V-�P�&�9�^o�)yLV=�mM��_�ccޤ, bؓ��!H�!���ܣ7�!-E��������t+��h;�x�iT���ۿo��9��"���~�G�����"4�J���8�/�e�٤x󷎬g	t�����pӅ2�uL��W�����>��h�X��G%�I������\���������h��	,���zi�t]���U�V^�]�2�F����KĚy����o�"�L(l����V	Q��=\��}�:��M$Q��ϼrk~�(t�faT��w%7��~pX�/h����n��5was���߷x���k,��G�5A���V��`a���
������=�B�-Ӑ\����{�5NO��"!a��po�׆c�ԇe�Y�z/Kŷ���?Is���CFt;1fﯝ5$��;�y
T~�¥�h��`���3����f�pNz/����y�ah�۠'N0]5�~-�lh��jo�(�"��2z���8�ȕ3�)�<��X?Rl3��jҦ#t�7a�H5�8*�ָA������V�-Q��;[A%�9�M�����Mls�_�U|�
������O��l�0�q�eN-v����Ȏ�@���.�����>�Vvo�*�����q��i.�Ȫif�\��b ����v�,N�4+����Yw�Zm5V)�a*䆆�Z��R!�[<�@�1���:���bV@�4N��hsb?�y��IEo�W4����F��:
Q�n���!�\�c��6� �-�Cvԩ�J���m�%otz�✓�2��dI��zXnՃ�p0�jD[=��Q�Iv�����1�˦ȉ�}�ݕ�䕮G_�![�rݘ�EE�p��)qai+LC�49�p��$��J�|(lv(��g�~��~(k�K�i�(�������?�E�	�W�=���7�Tn��u��o6{� ��2�q��������l�W�ן�����j3��|�8ߓa���p���E� ;6Ìe�.ì�X/2Ѥ���I�� �G�o�	���{]��3�tdF3�j�+�hd���F�AV+���.t�5dMc,���Uk[|��{���U�4dO���HO6�#N�,|��!��a]�F��TJ ��)C��)����vI�C���W cT@��3�t�Q)�(p'�h#��V�x�O�4�x�ۤ��;�-�H� ���qcN��r?�6��8���i\�v��LxS������2g�����w��߅&�K���O��J� ⏧��LT�+G�zZ�]k��	�W����Z�j�mw�.�T�$�*5�1(La�;��o�ơ��&����5qz65x�3˂b�$Wga��h�h�!�T���R�\wY�|�¼�
4G���`+��eN���֍M-����"g@�LY�&��*��q""�.��=@oX�[�J��~'�д���m�F����ߊ�w��H�c��O�?P�qT�mZF��	D��FR���f&ٗ��<H��!B���4�� ,Fa�w��� ��Q�h�"@�ԗ�2��c�����^��H�E�Y{J,�a����v_�WEbԜl�z=�}DvװO��S6�A�
�_���	z�r���~�ME�E����춃|�>��u�9P�if��G�[��)�>��54@b�y8�a�ӂ'�ژ�̏6ѥ�?�s-��h�n�Α�	��u��J�cG0Р ���&�]S�ҋ���[n�d��RD�+ɓN������o�ehWq�d��7K�)7�s5�*���\����7�0�@u/n��ć-�m��
T7�̎�z�^�@�f,��0@ ��Pn�&֙6��(ϴ��`��$&-
�K�s�g6��/ȃ�j�_���]E_�>gr
N�7��ɏu�4����Z�^ڟ��oX�l����L.��Ǒ�?"�bH���?[*��f�h���YR��5��uŧ���+��#'�|�T�Wp�>��-��ne�N���;_����$/��{ b��쉛[g����8��� ��
7�,>dt��֟;`������2(�x��X9z��%����ӑ����0h�D���Iqa�DP�#�z)����80պ,��'"o��*�b�R?&ZL��%4N�`���[�`��W�=Ʌ�A��ݶ^�Ow��CT��8��HO	F�����53Ւ��h7a�S,.*8~"���?�[̙Y�9����s��D�;� A3c��ִ�م@�4��������䟌�Պ�������f�aР�z�X+`����%:@���o8c��_-���ڇ���2�p�_�B]�/�L�$�:�w�|�����2��Uј��;�zy����5��)�믵j�5�K;^�f�hy��%�Ţ%m�������.���'�����N*�|[NY	8}FPw�Gw~� ���0J}���;��X�����Tcךoa��y~���/,/�QC���1���A\w����Y�h���p����ԊV��MB���=�w�����Xͤ���yAE�������&��������~�z���{f,�ŧ��v	�n��r�h��vSF�V��.�ɲ��C�ٙ㠔\"�b��D��)�ߴ��cHg��p�K�F귑q��ɯ�ų���������}�We2��RX�0y�n��m�u},�J�Zc�	�Kgޅ?:8X��}����3\����/#��R{�*<܇��U�.'Z�嶮Y"�D<z����Um(r}fZ���{N2� ��pR�^Pz�Ft�PX�.##y�P�?�`���q���\˰n"R�G�٭������M���ôhiq"sf����"����&��������hN3�������&軈s����/�z��r>�.a�u��!��J��F3NX��ȷKe����H�5�-0��ia5��|w�\7l}�?��q�R9FY�)?Iړ�c�Exm�Aof��C���i�P_�������S��R�wv�ΎQ `9��r?�����u	��.�����)�_m%���Uټ'qG���0\���&�%��rծ-,��=nXIq1�����hljHu��r�&1�L淸&�:�	�U��$LO&�kN��q6F:�wd�១���w1�<�e��&B�?m��g��cO�*��:�+�`L���H(L��:�I�i(e�˽���J
X/�k�(y囉�����U+��2���+ܾ�K�d���P&����/����J�CJ+�W�&c��)I��_��ў���3<�Zm�x��.%�"����uP#F�t�*����T8{�π�h���J~q^j�$2Y1�s��P�Q_A�k�l�	���33��B����n1�!� >���ɞ����}^�� -��ق����qy��4f�ש�?����IB�}2��<=��p>��|5|�ۑ�w��2O�_��o����M}
�[��?�L��;տ=V����1=3�nvt����}2	!����8��i��nx1�f���a�ZI�&��=��hp�>E�
H�/d���"�A�%셻���|ʓ]�km0�֓cde?����Ѐ���"�=aV��C�|���ٴ3[�#c���N1*�z;;!JV���L[4�4��e��dTd����-�t��o��N����U�s���|i��v�q�Y�-̧A�c|~�(ap��j�d�o�l�0�#"�b@��LaV���t_�L;����ٚ��Y�b�'.ww���.�5�
�Q}�5��ow������GF��^�}::�5�T���n�R������O��3Ё�l��m�SD�tn���ܗ2�s4�����^�U��EI^��3�gL'2�0�28<�X��PyƬ��nT�p�q�õw.7pDW��~L�����^��J��/�؜����P���� ,m����Z<��K�hL�q��q�������V؅��Ϩ��<I��C���!�Z��Ր�=J��@��5^�R��#&��X�n��|��v�5yG���԰O^�P��c�{����nga�D\�S\���آ�)�S)FҐ.4�CH�! 9Q�@��O��M�boiG�@��J��d��9�ߴ�,m�����,�M�"��V_���[텚���2D�>�N�Ƅ��m2�,�Ϊ�R�?܆�r��^r��>HA�)�{�-$�ڒ2C�1V	Jt�P��iL�'��/��_���y-�u�+)}�OR":5<��!gB�s���_� �9�jsƦ�M�1v���U^�emhQ���-=��9R9��ɸ ��6uJ��������~�
�<�*��b�t++ؕ���\˯�4>�%$�����W0��>��(N ��䥱�p�+�9�/�}�on-�,�)��խ�_ɩ�6)�*�%�:ZD�feɓ�o%I��˫&��@u�#�Vo+��6 ��X
�s����&
O��`բO~V�Y�0Փ�E��,$2��ЉS+f[��]�p����6�������֡�"���ۄ���W[�ѻ�6ܒz���o`
�����1r�@�!)�����G�������9"3q�~U��S��ʴ��3EdR�*g��R�m�K��ܴ'�@�Øpo�{(kgǋf��������_��#�F���̓5�1�5T��O_¼��k�������@�iHP��D�I;l�z_ �§���UA���8����*�k��)����v��kK�-X5��SU�����������!��w@Xb�<=��b�V���l��RL=l���v!w�z'��2�^�4	z��{N0��B�[Fl�8��(��s��LYnӃ]I1�xGAd�!�Y;ELn����䆥�$ٞa�lG:�@>R���t��G�#� ziġ���f��?�m"� l�יлv5+��v5̮��̶�ڎ͍.�O�'��_t�Y�����6�_7�����̐KA�6-���Z�6�"^Ʋw�8%���F7���/P��
�?fA�Y�ABoe�ŬjU<������Z�k�M����I5._~�&d�Aϼ�Y�},�p7��)c�Y�-���{D���:��+N�d*��x�O���X	{�p�����_�� �"xB�pɉ�?�**f�1f���Ȉ�������O]?S��R,�� ��@g����P 쯑�צ�õ�M�~�_,��t͊Yiy��� Fӷ�LW.�}~��w��Iz_��Z_Q�Ղi��F?r�3��u�J]N�
�|N9��F�
��$����(��������n�D�w���J�[��m�Z=7���I���AMpc�����W�;*a�p}�t5���V�c�9_H
'�#V�b��[W���L�ƚ��ybt�u���)pָ��l�줤o@�4>
9�Gjr�*Gsy��u]e/�B���&��	?q�/�2�X��t+va���q����2�l�ֵ�9�&a��D��+ѺA�}���P9�G$7���3�U�q�g.��]uy�uH�"p�ZE6 ����mϷS{��\&��'�����=.^�������]�P8��r��-����u�v���^�˽�BX�ၞ�G�"9_<���INq-xj����l��/pA�@Ai2�A]d��������odB|¹4n�.��쒮�k�	����΄��S�"�q!,���4�caHȇA��f~�d�T�*<G\��@*�h��˙�
�zʏ������|����K�O��-U��k�q�U3��u���p��g��+���f����ʉIRW7�+���0}�"�L�x���L�;�~8�?T�Ƌ�%֍hpJ%.�
l��-x؆���N�<v��k8oQf���3n��M�<@<�/>�8b,H�l7�3�=����R&��^n �hW&��"� �o�mR��y{�R4ig�a��8< �z��ȶ���ý���8�pO�P�eA5�J�N�,C����ܙ�Բ���^��`���T��҆307cr�ߵ=�ʢ�Cq���z��F�L.bR��s����_�h���2����$�_S��	���qHX4Y��'�%��H������:����_�ZB^Ǘ�κ�KS��:V��
�e�޹���]��;U�t���j<Iy�n�cE�q���>2�7��i�"� 6}��τ��'e�Ȕf"x�΁-��.�r�̡�*���|��V �&O����|P������q�r��͈*�ŠÈ3�B��{kE�-/_�yuD���!w��@7�\5TA�>1}mU��e�}��ݤE�@gǟ�]��v�1v�񯧠�.�q��FQQ�����S�@�2���W���*�2%�G�@549X�~Yn����J��DY���^o@t�,���ə�<ez�]N�Vi�ԣϻ�ĕ�x�x�y6%�.�%A����gSE�dt��u1�˗��w�S<*49�~f��#s�x�*�P�*��t^St�Ɩz3���v�:�c��ܧa'�ͽ)�[{����\|\e��t��Q���m�y޴���}�:�����P,�-Q���=Z}�>0U��z��Wߡ�m37(��BA���Jϑ�+�w���{+���t��aE����r�ޣn�؊��*-�;b*7���tѢ�M�;{DF0
�>Â�WT:�n���.�u��1�:�Wʩ�&�݈��!��\�֜� �~{�_�-B>jaA�S;�˳�'�ѽd12�k�K~��.�OD"����(T�z�Z����@eN)?\ٙ���;�'a���d��>"���]�)6Nq��X����̘dݻ�醳I��_���I[5۟�%�hT��yј��*�GW��������Yw��]�dA|H�a����Oƣ�Zh�y��w�W@�C �Z�ڧ�SIiF:�b|(=w��=��!x&�C���O��#�#u���w���\�?E�f�U���y��)�6������-��2�����'Fvی�����Cl����n�k����HP��u�ۈ]��g��R��>��Ӱ��)��[,��)x9�O3���)߫�F����H�����}O���ۀ���M(eN7�L&ɬ�ѳ��G-�L�P1�1��g���AUa ��J��{��+@6�J��u/.��ܗ,���,V���4R��O�Y\Fh���f|���6� 0�#E^���&r!�W]�4�p�T9�^�RG�~�>�W�k����X���J�˲Z��n�ȇ\>Ƨ�'h���D6W��װ�8��ܩ2�nB1%��G����H��]���g��F�q$Xr6�6�=���*ؤ)��$����~ �r��0�{��7<I�z�Z�v���g��U�H2�P�Ɣ�Ї�L��	���Om(��q[9Z�D��w�j��3]%rH��;�&5���q�YH@9=����+D~��`�}˿�I��d���Ӹ��k�ݰ�%Ź��裭01H�Hg��ξ"�m��!�f���~�����A����dx��]�5��������F:%�@ډ�J���|̃���IJǅ,��=蝄އm%H� �#�7�I1��is
�1��� ��<{=�B�"ȊƢN�Aɋ��g3�F�[B�Df�s��{IR_���b�D��K�V�����lQP�/�� d�iә}����[��;q�p��/�Y�uNQ��쪇��VT�;Qe��f��r]���;�X�<����qW���QD����̎�U�RMv*��˕\9c�h���������7lnރ$"���i�L��M�?W���Bv|i�O�
���0qr�2��RȆτB.�Ez��VV[����6*����Q߼Ȣ���f��Z��p*/S���R��`�-X�6?Q�{��k�NUt,�s�V;Qu)�/�1�<����j�w�lQ�>+4��D�zKj} �
�4!�#�8��\� �r7#��3��e����0(�,�^�(���mfU�!�C�1��)�K>���<1v.����F�
߯<��!�Ä^���/��1Iq>�5��~�f�ܱD�P� �w�8Ը3|��a�!_{+:Y���ߨ�~��R���?�(�[�����u۽!%��RdIj,L��v�@8Q
3�Dͯ�^�V�-����u��I_
ɕ��Oܬ���`!?��1W�^�э�ӚU�®)��ݸ��/��x����~�DPa����Ά��i|nt�����T���q�z���rk(S��8�(��	
ǰAH��mx��/���7][�ՠ��N����z^�EZ�{�^�#
.�I�%*���%�8�gw2}r<��\#�O����-�rШFb$&�HԄ՗�u�!L�'X�s����A������G��`��_�P��ƒ�Y�-���7S���py���/���� 6��,[9�~��'+\�I�\��l٭��g�D�p��Ǳ.�Þ*���q|/��p��"���wR�|t��,����n�7��n<)�9�*hΏ�ڡ#���>H]��tP�u���N$R9�S�vAb^TSl��4�ӰD��}˺%��d�\�p���׮��İ���=sC$��1`�kJ���H��u�t*�> U'[&��Պ�4��p�b7�4��:7��UA�e�?���n�Y<�rH��b���{:������=����*hPOY�zLM��믺p�v�L9�j���|����Q�I\)u��w�$%t7T��M(�*�ގ��1��(}��ej�'Vd_�i׀�"�����AM��@u�I4)���+������E� 	�.�cc�T$0�6�/V��s��Cw6����Y��৕eF��b�z��Qb����oP�$P_�*~T�+�5��ቁ��m6��6&?�N��lġ\�a��f�M��.�p �������4;�y<�D0�6>��S��/o�cSʎrWo|ae��-0n���;�Z9f���8�הc't���˿L��IV�X��2T��nhPMf�^c!Q��=�*����7u�q9X����<�J��ji�����b��4f�}i�� '�������i$�E�Q�;0�׺ZKC4��#��I�T����I_<�4��7uEU�I��l�k�]����v�q��ٽ���\Þ}���+�	��]�2*���PQv%b,BE�P�aah zo9�hw��� �I �,'`�H��;�,(G�k��z�a5lx�k��f���8�z��	���3&(v�����l[�I�nz�d>�	M��`1%٩�A=�.�v��+��>$wXb��MssR~"��R,Y&�'�,Q�t���ݧ4}	`Q����h*BLs��2^x��p2E������j.�V�e�<�+O��$w<0������,�����}�q�	��£̽������
[�� �9�L��]�Oq�-G*��ڱ�',Z�/�a^�6Ҭ�7�j�}�Y��e��IX���&HP����$�:Y뼶d�L�I���w��QAl2U���r0�C��e�!4�مB��J��%��B&Ԑ�?:GsT� b��_x�GM���V9���*U$��ْ�mAQ���g�B����]q`J��)�L�JI���'����6������[t������]�Kٌ�1}�NT�1�)�7ձ0m�V������~w��mK~a�I�+���ɏS���&�'9Q��+���5
�AM������~��9j �4M��"�+3H��("��,�/b�ڜDL����]�\��5�����;aj:#�p_����p�fi)Ǯ�GUڀ�J���;�����DY^֙x���v�d��D��x�^s# �r.���4Z�ǲ^^�9��N�+%�88~��|9�`�?,b��VÙS��b�2�π�����U2�� ?���B��dL8䧱v�����@	�@?��t:�e_�$�<5�\R����-�%$�ǻVk�ou%���s]�:ü�
��\�[�6�M�o47zmc����`3�19����g7���}{q��R����e^�QJ|��{E �U�H��+�>aın��E\m�WVߑ��1s����~�տ��ɴbu�qo�x�jEd��E�3Z�-�`�R�M&}�7�p
m6Ӡ��y�:~�!��+a�x)F
s,��es�; {�2��w&�9���Z�(�	�گxəjLe����yGGs(�!>(� �9?܄(�uz�����Kr$7!����`-����wZY��詸��My�=�����.��6��9�ߞ����>tT��Aw��.�+�y���υ�L��,�k��-3���L�qml�J�Y6�.�-ĳdz�sK��A����4/ ������f?m}c����f��v��[bE�*�#"4p|�g⯀mV3��n�\�Ãɝ�2l KuԻ\W�,�`�?�W���k�y���Q#��f˴5�6�Y��r�2.ⓌN��&z<��u��9S������Ԋ]\0��./f2�q��i��9-���-M9O�G����@A�U5y���A��	��՞)�AC�}��"���_x͠��Wf�Mt�#u�w�WF�����d3o)p��d�惈ۘ{�/�f�2�@J)A��K��'���=���Q9�\�Q]9�I���>6�.����ٳ�G�Dk����O5�M��~᢭4k#P�A���'��
Z�5j����ߏ�~Q��ِ�A��s�B��S�s	e�
�9�U�3,���yKVK~1�i¢��H���O'L�8��!N��z�z�V3aX�I-�$�4�F�#���c���5�)�>�7FT��b�H~���EH���-*�A<��k��fIشg�:�?3\�Z�R� XM]����W�U��~����nl�4U�6�A蚩��(�;��洆�������j���[n�l���	���n���m&\%��p�/�g�,�!��X�N�����%5�D���	�^�H䮗�,�Lh�}up��㑏?c�-]-�=2@�9�%�u�V��+�Hn��k�-PU�z9l�$�]kY���f*���ۺ�e��[��y(���7;h�+�dt�<�<��P����48[���;@"���Sxe[I��'��mB�\��^fH,�Wѽ�FP�L��A����K1-��t֜����~�R~�Y���n!X;�칁4x��'�F+w	����v��N_�7��sV	��XeŦ��*���(ܽ�T�-X:?�;��Cѷ3 6�etN�"Xv��S����ܽ�IQ��J:�r,y���#�}��9@>�?��RA8�u��o��c�����[z�o4J�D���.��Jai��z��7�xLu��z�&^3Y��0mg��&�m��m��t���'��q9�Q�E]���T֖���;Q������-j9�x�W�Q�2h���w�[�1��4��T"͝���|��S���
_�6G�R�+h 6]�P��"�@݆e@��S���u|��t&�1VD;���u�D��+�q �@�_���E4�/���T���b���f;Vz�����OH���g
mM�,�.�.Co��^j+S�IAX�s���#��MJ���}����?T��Vx�N�Nwq�t�V�/ف����n��F����uTE�	�z�zO��xE�fI�׆>���YsJW�(ֽ��)�s?�{�M�>v!Jc�s�����ZC}a������N���[���0�2dsַ!�J���]t���i�E�*%C*f2A���%��%�n�V��J&bw�9�+;���g08�P	�M�axZ���ޅ������[1tL�"�+��
�GD���p�#_ܮ���:�a@� ?Ùl�}w�׬ ͜�:6YI/��w����}c9X:�N`m���YA����IZ�����[SjZbRg1��>m�M��󗡔<��VT)r@�v�++2��e3�*��{����d�l�lM��)�6�%���5���[���&B�L�k�`��Ǖ��3A/�e�� �K�Y�J7�&C��_�a+��h �fR���JesK�J-	�$��J���1���g�-:tc�̫�{����C_oZ=O���Y��9;�ٮXEð�i�`�$����}��T�8u�#+>I�c���T�b
f�TM$BP �!D���苡k�4I���tszpu��n�f��3��Ʒ��R/N�4����
0[U�4u3�i����Js�QJ��-d8)J[h�"e�6:Zx}��o���P
Y0�bmȖy\h�
��RS95�ѤB	n:��T��b� 6��q(�f����@E�	�5]�#79���Ȫ\%�>3e^��{�^P�0�L�l���`�4���v#/�#��耻m9��4��?O��N��[:l+��6*�"�A79���Ō�[)�A�c�µ���b3`��� @O�vS����̒�A��QC�ޮ
JC�d�" M��-����yi-����|Pg�n�����En؟�ڗI����ٲ�*�$r�z(�*ynq�*&J-A"��1Hmք�:w�x<A��U,�+_�t6�	���y�Q�M���""��\˾W>N)�4���@Z*EF	��N���@��s���7K�c{��綯�WPF�R6��C�2�匲��'�^�Դ���֋Gd�F%	_�r8���g)���2�0�������u�)�T��T�����@��{�\��� �Q�ħB�ГV�c��:�S�?�?�������_��n�:���q) g*$%W�)O~g�8&�fq�DA�{�z�܇M~�h�
uY�����ǎ �.�f7G�V��]5��qe,�u:m���@�踕��0�H�2f1$�θ7�8f�3�j���-\�4[F��sl�:F��6>as�=en�k[��ff��-���g� ��F;�']�Bڛp� Q0V�� .9'��!*�� &Y;V����ϻ��N��ȉѕw���0�_�c�W��Y��O��#g�����k��>��#�p��|s�t��3O�|ym*��;�S�1#��P�<j2� (� �]��V2Z��.���y����d�	���X1}�)�i���e�׵.D�"*�Ƞ8�8�k������g�x� ��(Y�ܮ}�q�����e�~��T�W�? j�*T/]�:F��RbØ���
��I.�k���}�1#�����rx#��e�qG�vM����(�69��w�=\dp䡂�����C�*��yVS���p^�Z�����!^�\kk�!����gθ�7������}z��G�߃lsv�&G��p��b�� J2nT��$TJ��v�3 H�ԩ���_�
��v�d�IR�혶3�1��y��S_}�u��?k��J�ۉ��GQ�e�{�@�����\_w�G����/���e�V����,�d�5�B';gz��x��YR�m�s.�DE�?C�����Iᦖ>�Rye;���1����R��!�A`�%~�1C�S��0�j�������E��˨tŬb��������U\z.�f��򚿝\��f��̏��<#��i�4���ʞ%/�Qr(q�J�*�$�}/&D��I/�0����i�VM3�����f�_����"X�t�b�/Y�x�L��f7d��a�!N�T�xh�S$�O���c_�8��܃��)��i�n><ہ�i�`�ϩj�fX���1��(�Vכ��6�.DQ�~sO���%d]5i]HR�o(���P��SUp&h���(dB��v��5�m"�M����hn_�p�-!b	⻋�6�J�D�·o��B$-�s˦e�[?[WT|�,򏂁B�����Q;��IZ\�+������/�Z�d�e�+�4��`��i�G�w���n�Ab��nj�S��;N"�.�����o�x}�y%���5x�@��� �v���q��$
Z�����M T}��]�y��=���{X�F
^��1.��z��٩��\}�:�f��kVyű�J�q
��?nG�޵���wF�^!Wɂ���c >�iߪ��ܨ�|!�i��E�'�FZ���梖��[+���C/kOwC�P")�*��HY�(\b̗�GaٴPCEK8�:�6�s�:� L2��{\+XJyԅ��qu�p�_��Q�����C=De�Q�>n�;�d���0�Rc+]��V�Q���׭�v���������冗:vS ���m�M�p�Xv3�W�1/�OG�����e��B<2�)>��z�@^�*?Gl?���������<f�l�8��a!�m�/}���Iii@srSx��qR���_�Y����!6`P�+���H��ߜ��.�F���	W7��W9��+a����}B�O�G�m�@�����3�3�@�Ϊ^�:���)Q�1zmr�����ʟ���dja�4��43?���@Q���9�ѽ�,��\Z%a�@�5=�P�aM^R0��E��`���(�y���oWq���*m�C�r)h�n�z�*s_��jy#�]�uӰ?Q&I�*�X�(���IN��U��V:_w��§�DA�����5h 'o�` <N�{��F:j��=�)`�_1�Ӻ�1�u��[��e>@Zq2#~w/Y������,�:�V(8�.�6xs�҈O\�!�<����e ݋��R��%�q�%T9�-��ܳNhs#��m�Q�s�ml_YK��_�=1���}-�UӔ�'�X2H׾J���X8� A�.��DoÛ5u�6.���Y���޲oۧ1����?r����D�V3S{4eO0�5�p�r����M���d��Z�J�J����Zj�w	]�W�-��Leu9'N>:�,3B]g���W�]��qq���q���Ť"�=f~�3��!�k�bL�3��3P��eE���#E�Y�㋰�b�z�����/�g�j�jI�=������q?k��˴���	�?����|Pߨ1k|��ʢ��sOָ�0��+�O�7!��'��K�,D��F�.`D�\y������L�lq�p�c7+���{[=)��]��yf��� ��	[U/�Y�=7_����֖��Y(]�@_����v����NeI�Ns����h���sΐ��u��)��K�[���n�s,
C{�c3%ZW��6i%�[M]�al�J��I�:NjȪ�`C�A�/�>��V��֌��=��_d,O������_i�~���z_�`�"�kT1�|��N+��e:k)���_��0Y�Y��B�0�nCO�܊&�g(�h�>0ɬ��H��X�x��f(~��j�F��Y���4Z�/GUX8"��y�l��ֶE=���V#�V^.S�)������<�Ԙ��lA��5+�/n��l��t�i�����"~H�zB7�V���z��1�B���1:��ݸ�'�/g��v�n��M��6�b� /���-��U�nA��FS,���ϨiXɞZXQˎ8��k��G�Vμ%�EU˃��h)����WC�N ��k�t����RB�:6��U$��u�݅���ɉ����P�c3D�l��u��	OЃ=�DO��c_}����Ky/�y4����c�,ѕ�z��RF����c��ޑ�C:S`E�5��5;�X�L��ٲ��e�����w<@��n6�w�}ڴ3@�9��n��D�<�>�Ĳ1.f	�t(s��������r��h�0�����eA[`P�]Uw����gJ��t��3��,���vı
�KG��8�􃺻t&���m_� ��q�ƓM�_��,;�f:����-�!M��͚���/���3􍐼Ӳ���Ϝb<E�bgʡe��1���T�%���g�(p!7�i��O��p����Ul���J#�L�FG�x������Al�.Y�����Lj���+�8^H/��GK�U�N8�+%�1�%왚κ����yR-5�C���>8��OZ,�K6��]�C 4�.�
М>l@�O�sT�ٙ��Jט<�I�t����{�j�� b�-x?��Q���E�W�NXT/���	ej ;/���ױ��aD'�!���{V^���o����/��k��}���c�?�Ñ��͂]:|���xr��*@��7� N�d�3 �s�U�/��M�` �s�\�n,5�nB���Mՙl��,]�B���4z��n�}�뷇4(d���	(eO[��S����۞�dN3�:8�����0Y��x����ei�|�/���;c)�#3k�ĝ��kR��['�
����F����
�;�y�"�e���)�o�OO8Y1)���3*�@Zrx��Z�~qձpr �����:�5�3CS��ե�NU�Qum\S����|��@T�iP>��^KB�>C��|^׉U6ei��v��r�3 S`�_�"�/���e(����x���ݵT`6��=A�~RdX��B��|f�֡/�?��ߵ��̀Ɏ�4i��v8���$�}F���_��+�S�?���HXڿcE�W�����B��\~��En�|�H`���V���	���l�%z�)��A	?V�V�J�%UU�X|;��~s-V��q��ܼ����2է�P���p�z���{I,�m��٫�@��&����G��R\�����ʘɄ̓Y~����ù][x�?l�F2(���0���xusa��s�V���C`�<*0�wf��;�n�6K�)׬Բ�������q���U2�ӹ�ۉӇ2�C�w�R�{(N���d�[��X7;%1H9Բ����/υ��N���H�\Pג8��FA��A����JX9M��!�5��J�gg��e��U��x�͚�@�l�/靲�*�>���Ǎ#ܹom>�vë3��UE(ᱬ������� H����O��ĳƉ`5O�'�h\k��M]�`ХşAе���.qZ�W�͡^rH�^�먜�bFm(AO D�����-���b�-u�ym�S� �9�R�5�G���Fj�d{�n�����^=<�L+��3O��� �V�M��FƼ��R%8��	$
m���
[Y}NB�?�/AW��?@XI��-�Øy�עO��S�܌�|�^�kx>��Y����+�]�Z��յ�?(QQ�Q_�0��2�6+�'�I!��4_g+d�"e�i_7�l���$�&�m�`y:jΙ&J5�dƣ~�չxGVw�&T�U_b��'�?���L��������[c�m�taj��z��7v�QC>��F�3í�on��������ώj�?�3�>�o��z֨tBrsSx�.hJ (�����7��g)����m`}!�1�D��~tH��k,RD�r�����Lo�~ރz-&���k	n,!I�~�j:h�ү��i8+�*�q�w���!�_gTo�A@{|�/�x�73q�&�F�!�� J��J���F:���Ӈ�輂�kF�N�!}�Cч����J�r��;BY!4�_"���K;���
�L%�Tțn�f�Ch���Y^3S����C<����p���q^��
�=	2�F���/3�zg	��^�<ˤ�\{�q��J�ѫ.��|��Dj=I�u���RpE��W}3A���+�<Bk��:;��3�j���S��� �:�΅Y��$�ټ�X�`ʭ�v�����8��HE ��₆��[ ȗ����f�ˏ�E�^��fZӏ�I5���v�b?NK\m�YA����.�����yZ���\+A(4Ԗ\ZV;�HwF����}<W*�o�[�@����ā��)R�2c��6fk�\䰓�q�Cq)�ȵC��[�6�'#ꈝ��F���g5\\	���O|1��7Ri5L����N����Q��6F�_�`&�����̿6@ 5�;9X�� U�WK|r�M�E�!e����H����:	ñ�:-��,�a:�wq�I��#.#�Q��&eE�נkƢH#���i�͒U��#���Ia��*�U,_����!�0�m~]KR2�
����í���w��hw��oq�<�Wn�ȟ&ڽ7S\����0��N�#&�j��.�P�l�@�r�[�0/9�E48�`'���� �&ki�pt�*!��DZ)N��>�b��e̼#����q'�B�v�L��|�ųX���\q�]�c3��&�Nۈ�n�7�b�iŎ�)����?��gP��Q����E(
� ׁ�����N�!$�?P1T�ԑS =��❲���8aJ;�|����'�+'�C��S���m]K�J�g�4�����2�g��� �um��<�%�)�h%� �P"�v4���'P��9���iy0�e`EO��ܤ�mXg����ԆU@�Q�q&��
���z����h��������{��gq�x.�����(�$�UD`C�#�Vz����L��z��!�2pܹݵL��]U�@�ևr�`��EZ�p[�v�}i�1��~�?9k������֥
q����l#y��$$X]մb�`X�ߣ�
-�e����!���`����rT���{�<����w�D�p�{Y��A����Ze$�X������'���ˏ�}	}��g!���{�1��ࡵ��1��?�r�B�Ŵ��[,	Z���a�n)ʵ�/��}�q���u�h��-�	k�����1M�ՙ���۴�'qy�h��9p��u�S�C��P�$&l]�ȧ�o8�8��Wz��닐�8�);,iS x�VY������*�KjQJ?�QV��eQ�l՘Ǌ�N�����{�����7���"q%�M]��!̞	{�n�w�����̓��-]�w{[�u5��r�~���������z������9hg��&�?d�I��͚���b5�VM�w����D��'	D��C�*�Y�z)ϫ��G��OO�_�n���q�8�_FU���19^�F��!�!��V@e�3�YoW��g����MR^*�;����a�va�	�S��e߹��W������u6���(���E#�ݒa-p2�nps�|�m��"���R@����Sdy����6��:<@$��2x�������H����'����Ц��7��a����~�=���J�e��&M5R(�g��)qƐ>jR�ɋ�]�8>�����l2j����v�Ю뻋�co��M0r�x:^ ���! ߭n��u��)N�h2��@D騌H�Q���MO�3U��
(4�
�C��{*1��<3@���-�� �1)��sV<⟅v�l{n��a�%_�,�����rU/���L�u!
b��T�48�a�V&����.�Ó�V�
��O1;�<6�&��g��`4�N�L���%1��d�s*މ�9�	LCz��:��\>���C�5�<�P���m{~=ikObXؓ�v�_�fB�M��.��j9g���jsw6��-p�����W��.���=��F��y=�����8/ s�ٵ;��E�7���m��asP�V˲�;S���u���W3�]�*ӊ\ȶ 1@�LI���!������FQ��撈"�����[�'��d�m�5v-|����2��p�[�P��/��l~.��(�o]}P뾋������O�Ž_#۷�D ��w��%�ܩE�HEQ#���1>�g���������D9��֑vH��f��\·֩�;
�8��@�a>�ND��S;�èؤ8Ƭ�>1V�m�$4\�`tC��GGϥ������|�ɷ-�3��=^ps`��DHf[�]qE����Y�s��A��u�cS5Ūb��O����2]JdX��t�̟P�O��HlU�v6v����Yv-�LSw`(�Cv1��B
��Dwd�Y�c�M�H�Z����m���	�[��@�E;��@�EǼg���}�w�C��8(��y}o�m����#����z��,�2j�I���װ�=�1f����^S�+\�v �ϝPQG��hCN��_�p��uO�g����^��	�j4��ZԪ�Y���t8Q�s9>�Z�����b1}w�e\�/�}���ʖ�.����jg���%��:��S�E�c�*���!��K����ѰDi��\��N�	����&C$1ی��`q���kF��p��.�����Q�E�b�5O�^�r�p���+���t^�NoTO80�QƓ]��`�]����v+ޏ�w��@O���ϐV@TJ!�M44[xu�G����ez�M~o�o?Ϗv���	 4J\-��TR�J��O�v�ˋej����M�o�gD�(%G0r��V�S������� ȹ���M�L��<��s^��P,� G9H�8N��U����	��O2ƥla,d+bk�7s��[��lH��25s����)5ښ�/�T��Y��^M�;�l�@ӓ3�z2PH��jd��?�q�����OB9��@q:ٛQ������aW}��ZÓ3��}�N	��6��ъ���^u%���pR{���F4"��|������6S��+q*r!�d<��� �D2"ꑿ�~Q��ӊ7c�
I5��s�>��/K��q�Ӭev���Z8�bz61��k����f��(Ha��c�+�VjE��J~�.sIo��"F��=�����(iu�߇�X��WK��Mߋ�J�d ����!�����Vܗá���6����������z� �<��G�-:��SӺK�����O��tH�YΖB�P1����i�?xf�	��ȩ
�8�V"J��3���� �����g8**m���2F�S0E�1 ^�����Ř�ԟ<!����a1�0��G�ӝ�O�s���f�~PW۞���8�y�dP�Ն��n�x��
���+�M���_�\n�w��w��e.��פ�y]<5��y�fS��A�O�sV^#*�-dƼ�ϒ�+�H6�Cz~��m��T]_�nhĢ�0�3B>�i8zFTH&�l�HY�2�G���&���[��[Ǫ�X-��2	����l��iEmpd҉�WZ��L�Ĩ������f�/�<A�D6
�����	���v�
�y���U>���N��+��
�&зcұ5+,�](zD�.Pt�4�O|3���#�Y����۩@B����"<�4U�n����-��
e /X���w"���n�� I:��\�]��{0�{&�]SK"*������E0�T�@b&�ӂ��r��N�2�գ����lFl���嗃��h���'�6O�U@n�G�1�C\!38�	L����R�����a�7ޢT�M�Y�%#�j��>bݤ�K~>
ht�z�8?NT�/�>��N�H
����9?�[� #���w-����3d&��i�J�<V\��x�Xaƹ"��ѣ8�?�NK��!��UT$�9���Һoi���3q�g��0:}5 W^ύ6(�ܢ�P��D6�����#�Vg9������T� �#)�'���T�<"��R ��ߨ ��ĉ�|ǥˮs��*�X�_ͲJ�����+|{����#^we�jC���Ql�������̧Q�%��zOx��6�tӵ��34(�#|��a7a��?7I�|LӖ�w��r�-�%���Ia��u,�f�� ��$n�.}���g�IVoS� ������Η�zȃ��lѲO��.,T�X��|����Ɣ#]2��Jh(�M�sm��"�ȯg=u�-F�F'�b�FZ�}�ǩ���!d��lY�N��R�nV���������V>p�9u�f��I�f��')���Blž���'�"f���"�n�Ae�����\�7�E�L�#k�{��üe�W�H栎�̧ N	p8�Ͽ^?Uj^��>�^�ʘ׌oښ5&��)�n� �T��z�S�J�wS��'c7�-��l-L]��UY)�����3��,�^AA�����K�P��/���s���o�h�_@ ��.�F��-��I��{ۋ�ʬ��,e�<�&���o��}����4D, "��@��g��zZ���Ou�cȤ}��-�l�����ɗB�hZs7�.l����!�����vn|����[�&�;.R4D$uM����$���u((.�_�x�>�:S�Y�X�oie+��JTOY�M���g���L��κ�ץ�l�\�Q���ɕ���yߊ��&������
�f����@%Uo;ly�[�z����p^��~s�s��b��Q'B�	]+9��̔�?r�x����da�. M�K)��SW:����9��mq�_��d����Y��C�'"��o�����&�ڇ�{.����D=��Z/�3��i�թEW0_~=��@����#����uh�KS�<�)WҮ�m��ʎ0���V�8�e��WV�/olj��^iv-�Q�9yb���$؂��X�')�f�O�7�2.�MT�8Iƈ`T�9wYXA�P���Hq�(b�dδZ�u�O�hxc]�R1�N�:i�����W#H���??��m�2��[x�K��KA����r��߃ͧ°����i�ڇ���=��,J���`���RN��B��Y�/&� )�q����%�q���I�'�p5#�dN�"����!�՚5�>p
^��pײp�+Lt��t��1B�w�^@�y�?c"���e���}�4����Yk��M��¯��
���;E�V	!���yv$G)�S�`�;�.�_wW�oO�#�1*����@O�l�R�TX�,��GjҫP#�헳~M�'��T��u��&��2a��+���U�Y�^(��F��BC[����&I�`du���8УW�RmH?Gm��FF\]�w�ٯ�[��Y'����Q�a�V�b�:ۻ�g�`�!�厼�������ECt�������Q��b$$�/A�=2>�]k_>��A{C^U��Yi�5h��ס�e�=C�؜�ǐd1m۳����Z [���s��+�J�?��܅n'8�yN��n���c���rG���"�a�Hd�|?�l�R�yڕ�x�=q�W�[(�\> @�k���k��?�>0��.�s�D��'�ʵ:���W�$�OԆ�8i����\�UsscPZ��<îNEW`D���Q��=�<�ך/*	��N�r����t+E���#���V�-���>�\*�o*=Z�k_��HZ��6�%��BJOpb�	W��/K �=N���D�n�p�q�)'�Zu�r��c����8ش)�_櫃�D>��oR,��0)�dc5��a/�Y��A�,HkZ���VT�n�8WXB�F�C��I˭����֘��I�yT�����)/���N�VL�����{�q� ��p�\tQ(�J�dj۷ /N��d}zCc�ř�2۷|h`x�_���Sʶ�f�o= _g������;������l��'��xĊ�u1�c��yꧯ��pO+�T�����\�t�R���1����_�t�����"s,=Q���'g7:C��4A�q���*����~a9C���qD ���50�!-i�vK��ڒh^#�kw��]�ї�7_�.b(I��l/����r�f��g�XGY��R.��h+�DI]y�~ +�8q�{�y3�~�H*�@��Ѡ���^�wL@�(F �zF�z�m�jZ����H��ݟ�&O���ʹ�@u�4[	-Z��O� L+��rE�}��Y�>���ܔ��N颓[��/b%�[�IߡAjgD����������s��Na5�m�-.$�GzwOU���y�Y��ݳ��4��������hI��ݦ��k�e�G�"��O�������1���Gg.���va��m\Mϴ�g`I'1�r��Z�i^UV���U�wyU��"^�����ܩ��Im4z75���P��L����`c��>�0�J�b����aLZ��GNJR�4r:ۦ&���J�kPx�k�\!�a�|zQ�!�Ϲ���,�?��'Hx��gӴ�R�ޛ�b7-���.�̈́�NE��u<��M��D�n�<�iN�$F%��[Z�Q~I�M�ܬSni ��(3��)���wA��|���֌�of���,�;���]јŨn�I��� ��ƅj��Ɍ�V���3�jf�z���z��t�l@��t"aXp"B�g���׆��}�vV�� �ޠ�����6�3_�dĀ�B�؉������0�k���L梧�_�w*͝�����5� �[h�V����sN�Îǵ���#�==���������L��g�m|��O�ߕJ��(���Y�FR�n⾍+��?+X7��υ$ � (�@�{�������hqv����uQ�]��;ي�e�q�Z�[�N! �)r K�� ���t���|(����%�v��d1fj�&� ��W���%�j��z�şA~ܫ��-�����8Xj�����ǉ��c��zCZ���4:KuF(�NM�z/l�D&��U��{X�d'�۾�q��z��'��}�ӍR�̛a�{u�9LW�D��@A2��k��	�#�%0�'w���[L���],�1ɿL®f�>���'���LT~�Z7��(
Xȡ��Չ��f9d��V1��>|tB[���"DȲ�כx�͍�,cn�W�
F���T�[S�_#�|���-� #{�����{'�������X<�/T���y��#Ye
�v6�n�BS��B8ee��/8��%�y�U�o,��N����h��Y��Nrʥ@�X�V[�3�*��^�Dwp�6��N�8�L�J��#Au��?����\v_OQ�-P%'�����.��6�8���^��2���O�t}�;@H�6�4���q��OK~ݣʲ��. �#��7˼�����c8s`Վ��唥��#B��M ����($~�7�B���ً@Ƒ�?]��Y'��`6�;��ũK��L�	�X�٬k�_��	I$;�JδQpdCc�:�'��{�ܝ|����
7���	�ę�<ac�lX��-���1uTM�uWS�3�d[��.ǧ��X��1�֠ʋO�{	?ũȶ��Y���hUt�RF5��{��뉵��LA���|1��>ɛ�?�����C��T�j�U�����-Gbi^��\�o`!Oh��gw���s��P�U�v�����l/��o�o=���e
:X����h>C&@��}���e��.$�G�zz����t�5i���nK���X������^
)�}i-��_s}�:]6{�8��A*��2]���`xj5��*�狒��2&63Z�E�Z��2d�z%�iȨװ�L�wo�2����30?�lੵ9��Ͷ�`��<�mNr��#.���/x@L.�7�y8gd�V�y�]�M[�tX8���%�Z�Pxܷ����]�'����-'s����݃|�IR�M�B���~FY�����g�f#(�bz3v��:8iU����+�s�� c��|f����@[_����#l΁�D��6$?YW�/{Ԕ�N��,�������5kq��l�)��&�c�?�3h��A�J�N���岳������wF�4��*�xjq-�'����>�F� "=� p^N[�pc�P|jKE���z]=)�礈�
��x蓁R+j�&�y�Rn��\��r�Э��ҪP�k��l�$�2jX��ܱ�R����;����c�5R8�B�cQ�����*̳}�
y�Cۧ�}܁@�
��h	HH�b!k��B�
��,���I8����Q�o�mr%g�h����h#0��.e��x���떒��qs� ���o	�-���Z������n���OI�j��hu�$��h1�B��3+A�t�X`�6�P�J��&�H��,嶊?:&�{>-��6�	�� z���y��������=E���{���J[��6~�憾�� �ӵ�1�p�D��=fN�?����o4���v��T��ye���'8Q�:.�(z�~Y�~"�g����e��I�@b�v^�r�Z��`�l��K.z�q6��+�i���,h��B��S��S,��D|��~��o�b���]���� H��S�h?�h�v��	�k��E���̭�|*��P�0DՏ|A{�
��V�^|Ux��yU?�P[U�/���9�hu��unjR:"O}4A��'���ȡف0��>�9$�i�$�m��z��С��E��2��c�G7
|G��u�_��:yzݖ���	<��0��O �3\��<|�9|�-�آd��~{��N� @y�u���1F��v���{�Axka�������Be��a!�F^0u����h���re�N{�\���p'B�;|�̦��ֶp�����:MC��0���Mz���Q�x�J(���������]r��}�¿�%*�POb����A5s�/R���3PF�YN��;�UU��r�ǡ�ȥ���Y��lE+I�{a$$]�\1��(�������T̫�{�ap�%���;A�<_i�32y���˨��Mm;,��Z`,��,��	�o�����C�#��f\\J����ɩ��V|M P$��X�(%Xe�$���y�]�TǑ�f�d�j�$w8�s�ܸ��8��*	
O�,�_�^�2��R:�Pg8�л8y�r��.���t�c��B��r��Q���,)6tY����3J���^GT�\��{j!B����$�¤ Q]�bKs`�ɹ�p<�2�{���f�H�� � ���>�G�A�_0�cQ��lξ��yOP�ǋ���� �V�Rn�&@,��V<o��@������9+z�u��e^����F�[��,�+e�,qgg��d?��
-�Ys=hd��T����=DˉQJk	a�YmJ2��Fǒa/�`h���qS
����F�K@���j��Y���>DW����`d�YM��[U-�~q!1~EVv�=X"���RҗWt��k�K/�o]��h$��|��y�� �(��yZ���OuF�>�a�$^�i���0���?��dы(�*5��U�'y��n�h\7?d֏l-2����Ԯȿ@���ZP���0FdH~l�JUym�zUF�CE_(���:��B��t�bY��F�.���|�1��E�É�~4��&Y,կ(��kZ|��o�1GB <���{۰�HZ������w�h�bv�Q��qW��C~I�+s��LJJk�)]�}�,,�4)mS�0�F��)��Q�l4��c���@<�@�L�`�B�[p�0���
��z��~?�������S�)�5*pR>��鲒&����n�<��Z_}x(��[��
F�UG�X��$��?B�l\��n���}I��?�}�FqȪVtL�/�/8TJ����9?�rȺWp��=�!�c�����PuU7hL��&b=U��ľ���/�}>
2�A�������"�/���@��|��0٧�]��i.��*T_/����[j#����H�H+ý$���[�z��0�B�Q�b��l=H���c��3�]k�V�VaFn"���a���o�uh�80���0��fA�4%�
r�����ˌˑ�IYg� �&����.4�9D�/ڝ���
>G�:_�mXj�W᪊j*S��r�X�Տ����@Ƌ+���&cȊ,#*�N�F�C�9��JYѽ���ڹ�8ཞr4x�{g~ɒ$ �� �l權K��N�:r��~�28Ƅ�m�p�G��FX��@��*�z��i�_�dҭ�1{V�"����J�������&I�Y_�K�#�ſ}X��k��/�ÝϭD� ��]#,#�Q��0�,x_B=aǯ�f[e�}��= ����+�UFynH`�mX�(�w��>�\kiw(�Rg$��6X��5��v��w"P��TY7D���KP��s3$Z�Ѣ"�N�eU���w�W��Q��9
�#	�zrؓ kUX�Z�
Q�Ǒ"�ˉ_�����d����G_��6�oy'����Z<sI�\;�ts�"w��R	�� 9�
êe���.M4sf�d��i,D-(��cF��NΡX��HdY��z�T؍;�X���;��.�Z�)�:������y�$���#���|�HɎi�?wV�h����V�@�Ȍ5���ߌjX�r2�\5��y��2;eF+kc����z��2��s~)���P:Yd\��Sb�,T�� �J�$���P��p
�P
�#��w�E$cz?#۾�h��g^��%���4�[�=�.��N�R��M9;0[4O��I��6��������� ��%+3��xD��:������{�N�P(�7�__~' M7F�JNsGM�Tb��+���W��	ƣ�`����=1��E�
2C�U2>�7��?5�<�S��mP�A���Ro��Q�^�k�p�R�[i���P̵�����	Z]��:?�l[g���L��C^��aI� �������x�me�BGP�߈��`Ǻ���r9��,X3���|�J���<t�to]+�|�]�`r�cI�;�\6�6���b<3����D��QS�k&�m� ɔt�e)w*]�[�+���������zع�dqD���!�Ǒ]+_
<¿[��5`�s�Wh�3Y�B��m�R�� IGs�4Uo�R]�T9Wfxj��+Yv����o�c�?�v���Z�O���l�0������f�t�4+�,�
n>���8ᇿs�l�4O]W��(��ˁ���jӇE���ۿ_e���N���*
g��?i(�������|y.sN��#&0&^��F�2���sZg�����Љ-aW��a׌6��?ˈ���"���d1�U򏍘�HF��n���h��6���{��6�8�D�S�,`��G�؄l^{"�mt*��񆨆s�*�G��@0���V�?���Y؀Q4.$���N�|?|Gr�N����[Rޟ�ٙ_4/��#�$@�E���Z�?NM�����Bd�5R�_!��
�e��.]�+���=����5��O�'�/��ew�iގ�A'̀�h�!���������IhsN�ީ���j�|p��Z�0sj�K\�|��
͇GnP�1�$��V����H���eXL�-��PW^Cn�v���ހ�*dJ睆��HRA�A(�8u�Dj���4��\\����� ����@���6��/��\g8�����\�B.\�C��]���Qx�>܋E�&��g#�|�E����l�O�R��=�Li=0D]��_�2���G3_k�/I|0<�����"�8a��8�4ǂ6���_ V�;𒇅nY�o���p+�j��Ȓ�`yl�[�@>��m�;+��y��SP����l%����8�~�{�b%�JI ����6�_/ ��;��W���ˈ��N1��˰l`��/"Q�ܻδ|Iɦ�c��,
�����s��Ŵ'�3P��n�s��,��pJ]M�x�"�]�Ʋs
�'	�)��R�3r����@u�sW�S/��N��X^~�H�~jQF��:̰���EQH�ċ�0�xkK%���q��e���m�����ݹ7c,"g=C��&��Ճ��GUTz�ݼ4�o��{�l�?�	����暓$�>+������="�f�A&s�`���$�f�5���0��Ϙ~2\X�b �F95��F�X=���=�uX��I�X����˜d*U�8q�_+"����Ze�A��?B�E��,��
mZ�k���Fg�svC��(򲷹�tC5y���!?u���$Z�B��2t�9�}�n�rB�w=�H�+�����.7:Ie៨1~U��sN�՚ܖ�����1o[T���
����T���ط�ÝC��j��1
��1��9!~@��)}*S�9��zO�V_�MYn������^�W~K�k��uݺ��ISx6�s��r������"0�K(��փ���o������S�&��A[T�JN�fkH!ʿr�M�ݞm��:�n,���D<�X���U(�.��[�aY��1��K���ӭ���T-��Hþ��3"{�lT������&[R2���+	���-5�6?h�l����M�,��s������Amz��a����4z���|�]��U�B���_�;����:
-���i�,CB��aKI�[>"��-�K���`���/�l����<Z�!RUL����]��� |~�`���U��WF��۹�"���7����H����a��/s�{�ؠ2���Eν0*8_�J�8M8G�������I�����ΘUoz3�"m�1��`�7�]�xk��Qpe��b�[�^�,�IX
]������xm����0�zH�=�s�쵺�;'�����s�t��Y:��	7[ٴ����q�3/(c#�H���q|58��/�$�{�4�zA��/�.��:]����	�ц�k�Mu��X5t�a����+�ݳP�d'�y���
�cR\�L����B�����A�'J���#RA���8Ϡ8�ƇR8�k��:�,Bw�au�B�q�h.J,5�=����G(�k��^���xKhNՍ�2�W�!P�wPc(B�1Cn�+�4����5��Քc���yE4��%�={)i7���<�b���N��J������0��;`}��J�e���<�C�V�2��N͆!Ȅ1Oiy.ui�)����2.��a�l,p�?�ĮpDR`�Oߋ�w���x��mKb�,�zTd�<Զ����WC�b�k؟������S�eʈ�TsJ�����!B�w�6��c�i͟��U���o��A��`K�4C�	��x�a�X��"�&�\��D)v�ZS#��87�D��ܚ6��VN� �����瓩Ft_��_�Q�.��RD)������d�Gt^��,FÍa*�����T`n+���ã�����"�u�/X��F	���w�h��=�,.Z�=<K�)+�N�v���t�uO��Ǉ�y^~����-��*�A%(�I��9Wy�fɚ8�����Z2	���]uؐ���9נ�n�u��]��Y�����g��c���c��{��G����%���s�Z\�_o|94�2�?Ť!Vܗ��˂�5��mJB�x��w�>�����X��)9�E�7�1��H�еf�1L/���̡"?ə��K�G�8�@9��W՞�n�������N��ksZs�u�toT���+�>�o��2X������20���!�a�]�g���Hb"mo
$Ll#^.&7n�9����+�<%�p�Wa�릛kW�c�)^S�G�>�&���T/c�y8�	lw�Ģo�I�!�K7��zá�!,����zT҇��b�
�/���[y��w��A��'7���Q{��ճ�'�=dϑ}Q�*C>�#���RWnpu�}�A����ʎX�� ��܅=��j!�,|)n�,1�ہ/��&3`K��Q��<�UB~�Z�$��;�5F�0�pwi-��n��*x�Q �J��uH��9:w]=������+?� O�O<�m���� 	� r����T���Y_\oD��a����GB ��!�pf��],gLZzDΖd���R�����f�E���;Z����g`����ۻ��'M#�1�Z��k���)�nl�S� �0�mF�����BHC�I.kC��{%A#g���u�à��X����Q��Ey3��߸����f���H�$�v8@Иa�7��0I����O����[�лŚT;�\jR&�>���,�;��RT��R��j��GX��%��>���:�rM�d0���@��W�x5�]J�pj�0�C��o�b~���6O1Tԯ���=7x�G-c�O�)�^ě=�[4pI=-)�Q-d&4�fHA��d}��{�������`����ʋD�R*�7�3!������qސ��(5�6z�4�Xy1�Y|�|������^RA�_�B��jW��X� ���+%�FػQܴsQ�A��RL�D3�s�Tr���0\C*�$��Ľ�#�40�LZ���ٝ"���2�Gb���`�]��W��hp�bR����l��{@9�4�2!C�8Ɩ��nH\�%f��ҝX�OE��0�A��ϸ��;T�7iSA��d�	O���6����FM�Q��x�6NYA��JY�׾�xE�2^��Y��j��C�>Q}��p����p<��2��b�Tr��P�#g�L�U�9[	.N_d	T�t_����_Է-{R�}�B5n�}ϥ
���.�°�1��trD�����^Z�I!2K�2����r�E��`������!�l�ٚ�΢,�,F9�������6�L��$Ea�I����&TDs-�.�����n���c�4��	�eژ�V4��j��#1}2۳����QǨqU�Ux�n��I�1/s=�j���ݣ�c���晰���Ї]Y�{��a�ZDj��8L��ѺPh����t��)�?N����Oj�B�*_��GU;�|�f-�ۺ�Og�(�B�Rr-�&�QX:�N�1�A�K�P�c>R�H�}��z=�ȟ�If�nyZ*]��-,�GgDWw��ϛn�a��'�����&�c��>�I�Ih/��wp;du_[����HVx�Kn��f���,�DJT�ą9,?UM9}�7�f� #�n_öcUYtwR�(0	��-Ԍ��Ám�S�6�.#�񬼤D9?�0������z�p���:,�l�	���έ^��*|��$���L��`��XVK�,���A��JJe��T< ���d����Ќz�N�j�#��M|l�J5?4I����RZ��&�?Sю{�G:'bnh#ٻ��7q���ϐ�!"�I��~�E��s�����Jx�1t�/7�HDQ���@��ܞ��S�����w����f�n8����^��
�Xd�_����q8%�U�������.�y����Ni������yG)�F���-�{�mTa{ԡ qИ��Zzgeo�=:,T�$;&���z2O��,�l�b��p -��Y�:��;V%�d�b����%�*tBC�b���!]�䲰��;*��
��+a1ɲ�0a*`�򅬘��#_�t�SY��j���z�b0�e[�Nl�'4g1?ܤ��7��`��������.�;�GL�?��S*A�{$��fD����`�P��'��Z��5�O���p�l��ƪD������6-Q���U��A����3�����I����;b����N53�ͪO�A�r�B��Qylٌ3윸h`���&�Q�aP
B���9�k��k�Kd����.�J��>R��V���&��E��=��bx-�|�c<vFC]^"����,c!K���@T�J��06wPj=aV��1�,zbp��9\PV<��@INJ�픋ˌ����3�]Ⱥyl�B�廬m�ͷ�Q\z)R"�}�K�����y�+\Ŏ�g�\�E�)��i��0\'��A,&]L,���.��YOE�[ې͟��m�o���l*���7-�Ay	�q������n�>�����S�<A'�s+#}nY��UE')��c�����#Z2�l!{��D��1�1}�yR3�h(E5�#���yf��
Z7�}e�fY�����s��������d>-mu.�1�n�R��_���3s�Ԩ!�@�!B�_�ӹ�ge�����2ˬ�!��j�m#!��=���|I������kP1yx�)���o�u����x��q�ȹ���QA8<Q�7'�R�F��
�Ғ��-h:�w�S�\D3�� 6�"���⏮���3w�y����^n�$q�5���`a*6$R��:g6p���p/n�S��6c��,�a����������{�=�|��� �a�fi���;X2n����E
k��	WM��7^-B&�0�,̌�c3tZ��K0l#Զ@X���X�����xFs%��|8WY(eK�WwȨ��K���/�Z��C��,n1�������GF,.0
Z�Zx^d����i�c ��7�1z���z��M����=�!h�-�6�~D1�ɇ��~L�١�)�]>ڋ�[ਈ��W��Q��H{�7�G<���C))������Q�gNC6�<O��{�*pvw;����a��C�0=S`����mjz��';.����z��e��&�j�o�ӏ$�N��ܺ(Ӓjer�i�U(���
��?t2���T����P0%u)t,�Ջ���k�	�q�F,�OEW�r�E	<ij��K�۪?J�� �FjT%٠�{�+��P�H�̤0$��$������d��Y�#�(�B$6y�n��G�Z�CJnsu?� �m3Qm��3���H�p��ue�%��>IZ�������B�'�UM��эU�aO����6��{��`�ܰXy��"���t�1�7X��q#��.�@��y�叆�o@��Ћ�_{蔐�
�5����6��5�O��阖����J|�g f:+���U�2L����}���R� �/��T�m��$q�ȷ�z��� �n����/�a�	�vB;?�6J�"W|bX�g,e,U��� #�ڋ9P���kn7�VE�]ft��"P,ٜ�-1@^��-b��k�?:�z�X�M.ͮBM�>&�Pc :\_�f�޶��b�dU.�k��p�S6o�g��q����,��>�A��M����qZ��$p�I���Y���mu(n�����A�b���4�TJI~}�mF�j�=���F�ރEh6�c4/&<���B���fP�R0���=��yfL���7���%���d�oj9Gx���:!�����]�61r�L��ʱg[�l^�g����P�v������"�7���S�}����~L?���t�+�m$�nV��<,Qn���0��L�38�A�״���r $�6ُ�p��g���c\j�󯳝iTd� Y��d�(�D�[���ca�(x��B5�J�J5S�N[�c!��{��}�W2��a*Ʋ<��`�h�C���=�H�W٤�3�%%d�	]��j��<�����8����s��zp�d��$�Ý���/�7<Ǻ��ڿ冏$�o-�c�^��Q��&;3���L�F���ٺ�h�P, �&��U�:w��B7M!�'���h5�N�qhZ��@���YXQ��%pz�H�ǧ�d�?�M��/Ei��T�6� N�Ջ������-b&��_�W*׊�
��6A�O�l�{ΦcR4kL�`��>-�e��yz�̧�'!���k������.��A:�'��a��שd�,�$F�"/%�ryő4��YT
T��p�"ncrf�1�h�W�6�+!6܋vb��e������u�#JO�0^�|����1�Ngw�y����9�)��x"*\��)��ha/�`c۪/A��N����p��k4쌗s+HnB0`]��J�Ԙ�Y ����N���,W4R���ekNQ~��n��]q$���B+3�|��>9�<U\X���|qF֧��<s�|KlT�Xvf|���5�;�u-2��|U!;��Y�K�[*-ǭ�n�ݲ�e0�	Ht@����L�u(�B�.ri���@vH��C(w�k]�"?_~�+�s/n��ʤt'����s��&����LBZJ)�,��}�=�+術�_�砡^<b� ���N�VDb�?��<�:.�����>�_�,IVWY�����r�k���z�=����j���4���kݾ#�F�?7�|
����M��(��d0�>S���*����9����?�bp�WS�����0Yf�۬�g5Z_�\���E��1���ʶ��xʓ:��������h��/�;�sDh��ĊU�g>�oE8�z��j��Em�~���ԽM��)wgc���IG��Q��"�TY�j�%���
�_�K��%��`�hz���̗LZV���Y��/�$�� ��X�ZțI*Z=B��5 �d�,�b�R9�L"��F�B��Q*3ۗ��J��|��c�N�p�*�Y>O�8���n�bR��~�1Jy?t.$��-��ۗ���	.)z"�(��z�^�N�@���ߎ5�����TO��l	Hj����j;���fEK
b�}�@`-%B�%Ӛ!S'kŚ��9����þA�t!�����^r��
mO:�԰����6z��/� �V�D��H�O�C�}o�s�FZl"��t�	��HH7	/a����A�o:�8*"1�U��n�J��O�'޽����ץ��������oT	�9Dn���⣊1{vl��.��SW��mg�.�d\	
������2�&T^~����c��`�?s�a�S�J��`���ͪ�����1ũtD��E�L��~���B��~V� ?�o }����ő<�4d�ׅS���-q��̋Uڐ9
�1�	�Rmpx�DX��x&h�>y���Ѯʹ+
#P��/�-�)��N4�季1�=e$��v��("�q1�q��M�{w�W=��V�hƗ�b����s��]��)��74�0��Dj����c7\O'�`Z�Q��<�ӣ%ϼ �O�cUt8�J�J��=��&�����r57�5˞�.�`}���k0�v��k�wH;�M�ݨeϤidm]�-�%��R�Ϧ���z��t^6�^y7��#C�1�^��G7�b��M<d\����{P],H`�n��!1-�e����������ceԶ+s�j�U��ި��l�̹W�j#����8�/�'�,��j�ʖ���r�?��w���H���@ŏ��LYq�r5Xa������|��a�~UجY��cТ˼��Μ�������eHҽ%3���\���`��h4�A��\-$�A�v <R�K������.�C����k�l�����k�z����z;]��ЊQ���\N-:�P��X���wY�[�L�^��E���d��u���.��z��H��{����0<W7z����7����o�Q��z/�,q���Y����\.�DO=�!��w ��l9닭���p�RiS}�m����?�>�5�ƶ�U"ч~�=m2ǩ�H��8E��S����/mM;vF��I�;k��T�@"��dO�ĠRg:==�2"7%x����lX+���
Q�l����2��Z��T�*;�@�ё��Af*�J���n
�[^z���2#�&�V����d� ��gP�9��R�!��ˤx��Ǫ�������$���4�{��؞�r��-d���{͹ޔ�w����;�&��w�r^��Kv�� F�N��j����13���)/���W�[��G�nN�\9U��9��$(.w�%.m��K�AaR��?T�m�'���[�R�У���g[='<v�{�P���\��mG8��M�{X�����S�����%�9�T���wz4�X &3k(R[X_�\�!����L��D�Y�ÙP�6t����2)�ۿ�tى
�����Β3Ń�!�/�7����,�{ܐ�S;�����Ǉ;���rZ'�?���`M|�*U j���~ ��oW���4T����4�<��P�|��׎H�)��*�4z��)	qw�c1�PP�����C���ٜ�LF�:�Z��
K*��޿���ڨ�0���GJk=_�r��6�IZ*�t�A��7�"�e�(�)�Wi� ����pd����
������d�wT� ��y�n����m�l�P�ݩ���6c�<-�s_�&��{ v^J���D�.b��ꯤ#��D�[W�<e����n�r*���nϚՌ ��1U-��";�㝑����͕qn�,&��M@�%��L�JM��x):Ht�<	v�g,X����+��@�Ei�f~� ���pdy�	�T跋2]
'8~Ѥ	 �
~-"�U�x����I�f��4?J<b�� �<��}~�CU�E���!]����&5X��&�5��˷.�e����q9��g��irnp@��
��rڒ�{�p��9�ͧYɿh�ա�<���!)��F���H�kz<L����*q��@��ZCy����4�������ǫ#�F�4���(WI���-Û0*��{e>�j=u�(��CX�J�y&�쯭o�y��d�T��PTpa�E��S�T�L0_���;c�� *�<"�nv��}�2�DN���@ސ�{v�s��8���g!�����3Q�&���[<zj�0WC���g��#8gⓋ�׆�|�C*��ϯ0%�K!�ӎ"�)���b�\�������b�腌=�������ٶ\�}����uw��l��^ڃm�=����F%�������u�Ke�{V�q��������+�=j�EdC١�y�u��A"����ޱ��0%����Wk[i���7����ޏ5IZ��vp�9|�'0��*6
�}q��ޗ��o�4XǙ]��m�Y9�bs�|������ta�@��:��ŝ�ˏ���
Zg>}2���R�Z;���CSʶ���z��&�y���<S/��3༹��?�a�����{���,�$[�N?OB��B)�����Z�+���f`� ��:�[^��^z}����k�t4o�u"8��� �e�V��?��x2	b�?�*�V�v/]ԩ�����'���bAqs��2�31�	��rQ��>�����������x��&�S[�$Q-���=�/�A"�u�]qT�˟Ix�Y:@r�������wF��l}����ꭵAӞ��[�����T�}[������E��:��l��tň2���5��R}������<ETs�w]����s{)$}Ah��g�eT47/G|�+�Q��W:w=[�ف�3[T!��,���=��2^_n��L��z���"�pE�\3���:1��I,�Gw�-A��a������IHd:��C�sY%�7(m�#~S��c��Y~qb��
(��<^�@�7ؕ�A�v��n<j����t���B��JGo�P�����,�
��`]�\;�7�M%�C��$tҵ��6j�Y�Ẕ�m�;�"
�k`T�:q:�C�3��a�;Y.�D�ӱo6i�!��� C���
跁���i�L�^�Xz����q�긛�p"�44ը⑛+��6�/-n����vh�?�����WC���餲 �/�Ю�?d- 3@�f��]O���tS�*+��?��v@B���N?C��7�@�mh�p�.}꠲�`��lc1N�t�'��x+Z�Ը~�h\�5��Zoh����J�0{D4ǵ���UPs�ꙧ��Ĥ;]s��F9�ZG�=�����57����]�/C����d���D�w��}��ҕ!������9��g�(���kl�#TѨҔJ�o�p��;'�z�����Wr��d����6j�n����"�*���e��K�d�8����Aз��$1�-���}O�
�M��_��������H@�:w|@�UQ���F&����YC-kem�kWc�Ο9��D�D�r��{�>�!���-^�c�8�5H�x}�
=��P2q�b2&4��%ew$m�Jp81���E�Q�4�$�i�����m����"�n+��p9Ð�9�i�d{j`$�]���z8��ˏ�W�uɕ��gq:�`�;��܂l�MVM��m� 1�&>�o�s���j�V���!�6j��T�q�`di�?톓G���Q�Szh�b]L"p�{�H4n����
��^�fV~l.�BG.����Y]�I
�K^>���Ʀ��^~�s�ϫǡY�]�1�#���{�5҄
�Z0����l_H&h���ʵ�I���w�:ܮ'�=%�݌��̃XzF��Y)��NL"�_:f;S�0G�W�[�����J���? �^�u��>0**��K��Q��E�Hv}y>��c�0E��
׀L������%q��i�M�ah�Er:��.�i�����ǹ�����*�4����XC_�b 7�>��)� �1��6���"q[#�;bSF��Wݹ0�$t�����'�
	\v��}��=,�C;<��
V2@�a�Bw��<�7˶2"%�v2V��p����k��������8Ň��MJJ��Y �z�f��V]���W�8�Pl�.��!�N�Hi^ǩ9��Y�\a����)LP�p-��i��|��B����������$��΅��z��V���P:W���F�v�t���BC>� a5CH&��^��:��u7x�_�ъ�g�����l9d��S[f �frr7K&]�oJj%��֙��[j��F4E�1������O�u�����LX�Q�@��L�a���γSa�1��c@��S��̇^}����*�M<`Ȕ1o�#����D����?�Cۨ'��Ee�l�����,������!�:�R_���[��~u��$�z"�hgU�w�كI��K���UTܴw��n�qhݳ�g%AR��7O�����HKx�P������.�~l�z�T[hw+%3q4:��Ħ14���zܔk	MZP�EkbK��<�#ns�����z��7x@�sL�ss�e����Ǌ$<�6�N�iry)Hi(c4���t����Ҹ�`^�64	�IK��f3$�3G7l���<����R�O�=(9C�A)e�������IN�����#xP@�~���H��?l(F���z9�և'⺴�7���z�{~
Y�B��E��V�<@4� ��3���F��M���7s���~�lr����T�1������4�nr#`��� �����*xFpP��`l��MF�F���M���2_���0�Ҫ.������$ƘA����t�
Z�l�ʲĩ��+��hgNJ~RU�K,R�i��CM��F�m0}mK��ô)�c���E����e>k�0��!�Ēvz����l�q�e���5��oE���$v����p_�E�Y�_�*�rŊ�S�Ҋ�� Bk(5�̳cϱ�{Y6/m�8Cy�-Ư�&��`\�A�fc����u���v��vW��7&�m�1j�W��6�h�.*���L���X$� ���"p�a�̺)Rok���$� �3���10A%���V�c�l�	u��qƏ���KXc�]�	M���aP�t�nJg�,c�BGW�;���r|��)�>� �uyb!s"^�|�
ry5�/Z��.���������2y�k����������(��F<|�V�MȊ�3l�a������:�*=�,ِy���V�ýY���}ʇ�-��W�� ��h�j�N�kV��m��{���2L���c�q1�dl��"��H������HȄo{k}7�D�I|���I�G�F1� '�s����kH�T�,���������:���_�>��E9b���S����l�rUct-i�7e	M�W���-?�����w���uiE��=`w��A�Y��LnA��	T��sl�ܾ��S���(
�ԟ��3e��l��<x8���<i����\�F������vl�c]��Jۗvj��=���H_��H�������K�Gq�������M����|����ˤG�ڝ��M��ߔ��k]�!o�r>�ʕ����e�Cuig�z�x��>���Gߛ��$�N�����TG
Qx*ZR�����|0�+������I��+�4�󜯳D���)�A�p�+@�.ǅW߅��D?y�A�:H6�'�ɖn���/�1�-��-0��G���ֺ'*�F�RvլZ�pp^���!��| 36=�ػ��OރbԆ��?���$������?R�`��b�e]�3]����<�C!� ������ ��g��`��G�3ǎ��mulڬT��op�qSZ˼tR�s>b)R��2l�lJA�'��Ul�˦T,{Ď�ࣲ�e�6W`�c����i���:�h�T(B9�$�%�QC&�EmU���H)F����|��;��S��V���ܬ4�*?�3����cgŅV�=�$s��>���O�6f��)�A��B]Q�08Q$v!\���f@��v�XFE��h�eQُ=P��98�Z}���j�0X��|W�̗����ͽ�4�7H���1�FÚ2�)ؐtgq�6�H8��:T��Nc!fZ[{ꓻ�~PrI��W�K�o��)y�"Z�ׅ�;,�o��B�~�
���h\�:�y,
�Z1�,z@Fٹ3�������a�{Lai���å�|S�p-<>9�7U8��A�uX;�U�BiZ�KV�i<;U��#����+�Y��[9y,6�`��`rNT,.Ӏ��*��'�f��D�����9 R7���6���0?o}���ZL�������@����P�A�E����R!��&~YR���n@1����y�5���٦߰�G���Eg�
�U#A{�ذ�W�N'��Ks��5�����'��k���t#�P�� �y2���*�;
E�]^L�$<��`��z�Ɓ��䤔n羨��ʙ.;Y�Ţ�(�R"�D^qF�F�9p�<m^�x������ᶚ�&��e�]�r;���O�D��&/{�2�����C�fvbX�R����	�!������	ǟ�ZMBA�_T΢u�9hr3G}�gĢ^��9�4�����x�w)�25�W@���]�^�zYv%�q�k��5��M�v:�M�i���M(~P�{<�,�T$�h�k�7�'�����$�|�c]�O$�|�V����Ft3��N
�\!G�n��r-�ҫ݌Tت�= ��)8�:Vf#9;Ƥ�Lҹ6C�
KGi11&��1�O\��w%����2E��YB[���M�ci��A��k^'Avx0P�,��lV*Sk�.��{�"�W2x�Z�)E��Q��Zn]�I������2��CH���)�>�%Z�{�̄���^`rK �H~�'��(v�ɟ�,.w�����*Y�Sm��߯���B^��*vv�|)�Fhp���#�R�V�a��y[�֧�qK�V]���䊵�}#��@�ȼk�6�>�v�,��]�������Ն��T�V)��j�p[�y`S9a��L(�Tey��X�v%�}��WU/i\�x2�$��������Rj�����^��}�yjL�f��l+���	��%��C6U�Z�ā>.�#^>���ɴOGT9$ɖ��j���ٙSꪹx�&zU�lL=`O�2R?X�+�Q�տ赳Gi�v����٧�7d�4Fn�xz$�h��w�IVЙ��=�� ]&����"�?6H8���h<�G�u>�����qۅ{�C��ŽWY8����ܳde=+CNqO��$+V��iX4� ۍG��H��bmw"��A=#t�h̽yC�GF`��(Q}��|�y&4Ф���E�BtuP%���QB���R8V6�^��	��m���y	�l��=��6�z�T>��"8ro$[���䟪8.c�2O�TU�(ӭU�X���$�����9� ���ܥz.1<~eJ�%Y���,jr���2E~��OܴbA��l�r�����1H�R�Ɏ���-vD�Y�%u����2�N�u~�k6A��.u�<�]t"���3��E��d�瘺Wǀ �!6�t��Q	�'7�Ƣ^���Q\��<$يS�B�>V ��;_���Xx;v��V��7E Ah�!^�H]�j�Au��t~�T�T��S������x.�W��f&&͕���E���z���T�x��4���v�BS��4O�}�������w��(23��a��8���푞(�t6�y�޺�0�{��b�Yn��b�X��,�1����;&�,V�3����d�1�܆��f5w�|]ԯ�������o�m��Z��lJ�װ����n�^����y+Bl-��j�/�{�/��)[�;����ZJ��P�pk	�ِ�~�,�.lҷ�?>W�~��e�r�	�]�/�b�W�"��a�i��a]�:�����ޕ�oNr���\�s9?�XV���i�� M�{!�t,�_l���'Dq2"����O&��w��$<?:��Z8�+җS_*y��K��/������ �w�O���)�zl�75���Cu�]����WZ�&5�V�pM�ms�-EH�~�@ �z���2��"��y8~Z�Kw<&��͝���W�M6��,MT=�C�Ta��א� ��T�I�#��ze�Ĳ�����p��5|�cX1LTX�Z;
}���&�q�X�Τ3y��?{��w|8������6��e�
Su0��Ƶ�&ň�*�J1�\$�fո�FMN(��/@�z�<`�>,�C�u��&�8��W�k����bo�� �����;ͮYt��~M�z���5aI<99�aY�n�RM��T���S-pqYP*�"y1��g�=IW�����EL����["7�P"�R��bSnk`������<H�,�wt6�+�7��F�N�<�®��W�G�ȅL�^v��>hWKσ)��p��i2�#�Gj!�|C^hZ�'ʈ=D2���8X=7�}I��DKT��:ͷc������0v�p��p��,: �8T��*�`��E��� ��ӂ�Ad�۬��$ǧ�s٥l�X(ȍ�F��b���v6�_U$nB����"%�7��6�i}����-����/�c�Q��8?u�D�R�����d� ��{�Rq��� �`a�]s�?*?��g�4qW��#�I�-�+�b�P����]�LD�U�!ܯ�	��'֢tҿ޳��	h Bq(�-7L��i!)��N�MX����IqD>&���Y�q���@t���*#@C�E�]wW/�'Mt/��1����'C��zbF��ß�:@DW��j69�����%z�7��3�z�x��:4�j�<״���*����kX�L�#�Ҫ~�aܩF�v�ɆS�W����q���[��zkӚV��|V�3�R�/wC�nI�.�p<E�8��zб_��5w6�ɑ�z�~����qQ��D/̀�<�y\H� ��
a\�<ͣs}қ��8.�(|�tO�]���Ҽ������V`��.�Ty?�����+m֯� b%ָ��O1h綁�e_U��v�����ͦ��(�����>Y����c;����U�C�d�z��X��6IG��=Ѯ��|��#�$D�%���ϖ�W��6`�Vb��(Q�� JJ7�wi���'^�{��N�-��B�W�X�ym�:��cH�d,g-9�)�i�`�#޶VB��_tѰ�X|�j�sB= �����C�h��:��(���Z��GId�%g�ͦ�v=JC�;�f���6-.��î�b1��ab��-�=,-Tpm�Ԃ���FoT�:7<Oo\��j+ut��D/�ІQ}�6yGfM@�]z}I�ڛ����&zԳ�>�A�!;�+��^`�9�tF,����^Lvr
��\K�� \QPHWM;[������a���c�[ݒ�(��"kД�"(H�Z����>�#0��U:hq7�{�7��5 23�	QϏ��f��"={�Ty�7�� ���3~���-�?D)l>3�Ɋ��]I����m������CjBfO'�?�h�Z�Ȱ1�S[����"���Q�@8O��B��� ȣ�2��we��:M�#ⴄ�r�h�?���o�p����񶋦U��X1�$�[�#6�I������u�f�񟘉)_a�"���Q��IڵKxn��S�P��3�������ov��?:OJ��^�8�����{�����{ɺq�,Cm:�'��kk��K�gA2z�y�IP�����M_jTF5/^fTۚ9�ᖓ`�E�9�<s���M���::��bs-��ª��i7���W�_t?N���z�L^��r\�=G����M>eJq��N0	i;�=��gg���)0�D��|knF�{��Xn}N&T,^���a<q�Ej	�G��H	_��m
��h������l���*�6|@��P��jg�ߴ�6��'Kn:��L��4�i����]v؃�����,�1*5�._�:�B�^�!��^�;i�(�[,��)񓋖Ɖ�����*�����"Ӕu�q,P��o�;��r�W1���������1�v���%��l�� �.d[������ݮdC��e�`k���GN�,>��4gw�ȸ�=Y������WoI{K�b9�+A�J"�x�D���y89Fo�NT���[:�=_�����ޥ��l<�ə���'���g[�xl�7L/<0�I~w �)�����]UD��)p�Gȿg��Ŝ1�fb���D�(@�@m�?@oV=�.�����^�����AG��nAȻ9�^~U	������L���ꏿ����M[S N������0��*�^{W��d�Τ��y����i���[�쾲blN�0��4���l��&�Avy\��`�O��-c
��o��S�	�˃c��ڦ�����2�����ܰ��M�R$R-)��q�G��P~�����Ҟ�O��H޴.~���]�1�7�����E =�6'�j	���wѨ��1�E��>~�c�� �0�3Zw����	׉�&�\i�����������7�xI3]4�.��0��ِ����Ώю倵k>�I5�=����9xe�.S��er8��x���y�H���0d���%�!e��?I.�^嗑��&J�WJ�: �_]ϫ3��?^>�H���91�
J����9+�7�5����{X,��ɀ���P�UH�S����;?�����bg4^M&7\'��5`1� YT�Ml�=�g(g9C~� ���J�Vbq@�*n���tQ����a�����X&K��ٌ�%F3�͔�C���su���ݴ�.�2q������!����sYص�}�ڕ ��q�u�=��\�\(��@�׻T5b���	p�`Q;]f�3�5	#߮͔��z��P!�S���k�fV��)M|8��a��{���������q���O��Q������A���5w{���R�M!]�-V�xL� (q�	
�Ѥ���� l��, �Ix�Hc�b�QК�?X�l�B$_2��ݯ�&t�խ�����������$+��Nry�?qʈڦ���I\15���A���g��5�<I�N��1+�\��K���>�W4SI�\��|�%*���	� 3�V��Xӹ7c��!�
C�J��je�d��.�4P��N��Mb^W�{�;s�k�s�?�e�df�|�蠝���I{��^�ܺ!��a�[D�]���Q��υ�{I޻��� �ϤK��(�(�j��(��T������[���r0�N��j s
o`؉�k:%(��"������<�����qv��P}�x�R�4D�&�؊�ds2�i�i�S���]�1�\?�j�M�Z]�G�[+�M3)��yFв��K�W�2fƅ`R���I��P�I��ٔ{նL�(e�'�D��������|���:��t�nHq�n�K�fU>��n&�%o�-���W��o06%S�b�p+f�[`��Q����c�DX[����!,�Г��m�h�;b�������q^��P����&�y�|?�&u���|m�g�,6�sp;t=�ޓ�H�"�񝧡����a@s��P��G�(��������0C#�$�<l�[�w���7;��v��/�@�B]��4�c",
A��";o�t�t#�|�L��8.��2H�FUٖB���d�{��)$2����H�w����f�,��Z���wB4ܶ����#S���RH��_@?�O M�Rm�N�J�������߿+��j�g�~[��-ců⹺2H.��d�9i{��p,�3ts@c�T	�p '+�W��%��~�ʊ�-7��<oӕ�0�:)22%Q��ì	���\<[�!�'� ;29�b�S�P�m��}�a�ʤ�L�����gl�4��n� }�ɄB�NF���}�̖�
�f�p1}��M���^�h���xzd� o���?1��4T� e�8��ƅ+�:O���p����¹Bq�"�����Y�=Y�ȹ,%��z�X��~���ڒz��n�h��, ��a0���#�2��.��ii:��'aǔ�sA�ӧ�y%O��I����?`AF�p�{?RO�m�����mN����G�W�_O>�T?��#�n���ܽ�^p����l3�1w��:Q;�s+0SeR�E��+�Y{��q�"���$ Fُ@���y0JN�~^��	U���p��o�Nd��Tvq�K��_��/y��U��&���6�q�tm���m���/)k1��W���9Gu��,%_S4�?�U���{��g$��s�4����YpA�l�L����J�a�%;�OI�H�ǀE"9U��_ӎХ�����Z|7>;�I���#C5܉����@V��]�o�"}'�a���y�����u���� �禐0�c�G���9LF�5?�O�,A�Y)�^xSko��m�CV)~�+�&&:�3�������.���H�t���H�o�K���%A�����'6��¯a�,Wr�_$�.B�͡ph�E�hf��C�Nej��j��]�&��G�{�r�/ű�`r&���Q�
��0Y�1�IL�o^4Y�R���5��a��
}콀��~c�!iVne�Z�@s,}�Sۀ-�0��������x]�?�rB�ZZ�٨�H� �ei����RUAg�	}q��r����.�5uԎC�e����2"ʇ�_jPQx�#m?]�.et�u0�@t=8�]lP���\xU���{�9[&��Xv�(�9�[�� �����`��H&����������ý�A市vt4��~�~��Rб漸��U�[=�3�rHm0�a���?����L�/�SS<����і�m��U|x)��k�� j���ѫ�:nX�ii7�)�LU����b6��s�<�W����&B�b����2N�i��h��\��e&\�b^��ֈOI2?L?c�m��?`e�|�$�b7w�>�po�Tf}ق@M��n�=z.��=��@�1h�~oڜ�9u2�xM�m���vʗ1�˙��ʠn�����*\��u�8#����������ǵ}X��<̾����?�F���&)�X�O�cQ��^)�����i\4$7�r�2�*�@5�K��yf�>�
�>��"�B���p����������+]������T�`^���������
 Z=�ۣ����Ά�7t���t�)0�G7������gCDҁlӠK��y���u=�mNӥ����+���̎�)�~[%S�����YΌK��nV��U^��F�Z<l�QX7�z��A����c��#Lg�l�.^�(C$v�oO2�k�|��q��8�XL�������]1����/��\����*�*}Һ��>��G�-���=�qLчE]���D&�|�I��Y�T���I��4i�9�X1�U�c�0�̞�T��|{�~��cC4�gh읽}�})+�P���\~=���	z1@����E�R �0���8�c��vC&@QN$}r��;�W��yD[�c`pK����.��*@
wjnVx��l`�7��y�89-�l�l��۰r�Gօ	f�WS��V�]�j���xс��b7������eh��qֵ����&p�]�	[f 9�p�]�-c|R�CC��?�t��@����}��iy*;���8�N�xJ�9Ҁ#��)��<D�EmZeW�}��߉7���=�T��z�R�A�>N����{=2
+Z�!&m��� >�&�. F��sqF�=y��l�OX��z,*��7@fwӖYB�n�?/@�|�"��1�Go�A�E*@Ѫ���{F�����l������Ot��S�74۩;\�B�	hE�3���~��)}4⒑����@��ɹJ2lE|�O��l��h�ӓV`����Y�2%�-7�mʭ�d�@"�7AB�w�}DB��� �vW{_#$�[[N��LKD�BJ��7ޞ�X����to��w
a%�	RtGe�=L�HrZ���H�B�gF�
�؂�\�\KU^����_YU�i�Ò�3ȷW*��/ZM�,��93�v�q�8��J)O��Q�}}��\��f�Y����[>f�ȑ�W~���I홮�D�w�0N9����w�}؍�[V �gLgD�p������s�8"w�	u39�ʳȾ��-��'�;�[��~�E���g}|�=�^P��2�y��WA����&S�rtw � sn��l�ʡ������|f������;Q�ަ���,��^GX��)T*<������4��(܈�Bokh���a7��D��Y���=�:�S%��Ҁ��B�ae��S`Ty������#��*�f�ⓚ�́���8����"}>�-��C� {ʦd����=��X���1����F4@�W�nEbY ���cr&;bK��3d:R/���/�M't��!�p�`��?e%�-�s�F�����{���V�����K��ޫ�R(!�Wy� ���	k*�Na�t��?�=zUB+�iIR<���~��lz��y�u� ����ߖ��q�
:�th� T>�@����
��\��3d�UX�2~�`ɩyP����I��Ը��E�L;D[eF��OH�w;���t��]�y%�ï4��\�3�t��d:�J�+o`����!��%43z��
@z�WM����7a=[�. "�<9�a��r�u�#W�Վ3�tؿ�A��|/ѿ^��>ڢu�&�&����+$ RW�slfn �O�.������V{[�R�ȯ�L�ϒ�G�d��\�4��8��qkK��n��,aW�K��;���.!ƂS@-�Z4y�� x����ι���F�y�~�����2����[��a3^��������l?|S[�#J��G�B�� �?���h���F6PR����S�*���1�3�*5��l�C|bq�ab1���!%���pi.���w&�p�v9�·\�����'�8��+B�o��OG|&Z;�"&�IiB����<�r2�f��MՒ��k#��H�㈷�d��x�RD`>7�N� wI=i�7c^H&8(C��@�\�u�9��>�G��aCD����I��XF�T�q�����]2<�pF�����9�����Qk'FY=>ũ���\��G�-��{k%�P��M�Vk�[�}���ck!j���qNx��?�9�Mi�r�LzXp���\%
�<>��OA�J;�JZ�8{̅4�*����kz��U�=u����i�V�hlzǒ�3���;�Zy��z=Y�c>�,����)��!xi�*w�A5��W`;���� ����OZ��Gҥj�w��7�Ds�v�^�����0��������P��Esc��4<G�5��6"��<9���b��!�j��hn�����7!�y����|���3=���4u��A
�e 8y]z�'c�<޲S3� 4��в-	ޛ�"e��~�g*�]!�kٺ{f��P�K�Ӻ�!��u�FN�I����������0���ׁsĆ^t{|r;i��_���B��v'��-D���0��+��Zr���OCq����Ԡ�>�G���p�U���[Ǻx�C���7�?@�'�<�@M=R��Xu�C���z}��r�yX��v_�/�7u�$�I*�Vc\+>A�v���c	���V|��Er��Ma���b ܝ���sH`F�;���1��;]�p�@'T��~S�qd�lI�sy�d������W> ���D+��X�43鄏L�z�䉁��kH��.y�� �c�&��{���xY�d�^�|�a�0oʷ����d�
��eN\����qpv�&��2tV�3�9�'.yy,�4�5%T_�����p*!@�5�$��HPr��%��m}���Z��_��j"��ꪯ�j�NGjmIi�l�������Q�=��ֹ�af,�gAL� �m~ӆ�����b���v�K�؎�J��H�m�ҥt���� p`f;�g:cU��j��ͦ��Yt-/�:�7����s�8R�� @�Cf����铺�]Zl�!2����:?Q�tpޟ�_��¯+t�ۂ����گ�'��X�i#�ڠA�&-���Olr���(�[�h�l�0�9�D�Oo���(è�eX�����0���2�
��/�t��X%��s�:��^�c8��i���*z�������,���_���7���vU��K�iڡQc۵�\�I�AC�9�����X?��'�8�g4�H\�>�pa�����3o"���)�.�*���E.ĶH� ��ނ/��I�5�sΕ�7 {��0-���.I�[��H�a�8�����
xn l�{�T^%�mt�t�B��Ĥ�����`?�Vp]7]m5 Hk�=������/�H�+jm�5��?+�׌��F�Y˱�o6�]��}5�4�s>���UeX2oJ/h2��;ah~�S�KE��uF7���&�=�����1rL�
f���p��"|f���l�N����;?.��;�.�P�g˒l�;�2���c��b$|L�X�D�/�W�#��Ʀ�������'܅G���&�oh���N�A
Td��a���V�*0��V`�@��b�}�N��x��đ՗\�~�ۯ_h�Ì���y�ΚFf��l��*�j�L��%�9M��\�R�+�ѭ��mDs��gh_�jRӭ2�z=V��ǒ� &}��7c�+�f���K94+�-�X0��򥯃���7��ܰ+�џ��|Y����r�gt���t +9[i�w�*�$P��t�(��ӻ�GSd�P���`������E��p�F�`��X�D8�as�~�h ;\}˚>�����'!rө|�(V&��g@Y~Q�1�%Vğn����8����2R?˃��Hq��Մ�����a$�i����p�"}�p�L�;�Y2��E�?��W.k�d�ܶ� V�+�n`^a��-����K:@����W���C�?����W���`���"4|���O)`{qGҸ�y��&{x��&l�̣6Gl|�����H8��]9�#�(�CQ��"6
9ܬ\�E��q,���Se`p�R�%������t;��q����OY��y�tC��>;�^��� �z�հ��Xc��i(�P(�K��Un���m��bo������z�v��	ٖ{_�hrS]��`��X�K;q�_v�\aX�b�٦���<�_eS��3�\�c���v�<��]+5b|�B�(��N�L��=9�ϨC�E,��6č}���uQ��iIdێJ^#�-LrҞ�_���1��="�O��|%�Т%-�D��1ȇHA���D�.E�y8�@����p���?e��@r�թ8đ�o���0���e��ϋ�G0n�3H�]e���6s�k�h��G��42³�1��X-��.�Xm�π�j�� 1�j2�n���(�o$�����Un(����C�Q�c�Y0�|)�jơ�^��z��놆�lU�Q���1���W���O�o1���':N3p��I&	��%ޙc���I <�î�b���f%�"�vbB|<`�;�}қ�m��#㼲�Ga�L�B�G�mZw����qǢ\`��c��ES>�k��Yl^ +Y<��mpP����н�&r��,P`赥+e
�Iⴽ�v���]!$l�����}�\�'�X_�ػ�3���M5�?:XB'b5c��u|�q�W(�R�DE�+�5���ˈ�e([��s�ݯ_����N����z*���������8�G?R?�D%#yL��Ӟ���G��Q��&B�!B��}5�"�����*5�a�'�=K4�z��g�+�hWх��Ĥ}㐙Gr�lzZ3x;��'^��Gp�[���Zvw�yX� Ʀ�E)Bs��P�+ϩ���!]�A6�t�����7�������hx���1��T7=!w�b���a��������Ǳ!C�棽���%��.O��K�����n�����w@�<%z��������_)����K� s�]����?��|��� �_ؽ$�F(T5�������fȲ�)�0�Rǡ�G�W�#�n=��iDc�t]!k;aߞFuQ7�l�L��"nd��vc�d@�43eZ��O�LGU�{��Ѭxwk�������se.-T-�KńO�B|�J�8�AhJ>�a<�������^�W���	Դ�N��3A8���@
y�|_$ѭ��<��m�R ��䐱��6�Ø�����Y��������P)�EK�0܉����}t����s'�w\&7\�X9�1��I�FF�i��>�����9���)[%�ssC����l��IQA:�\�GA?���2NsGr�;8k���$�چn�FN^@+����=<�e���aG���-X<�#�}Z<�4_��z���	��%y6��.����.�k��3� 
�s�^Ʋ{].��=�8L���T��Y��:��e�y�>W�;��{���^(��q�'jB�H'�`���.u�E�# !еґ2� ׷�`�֡��:/Ǽ� 4��1�5�+�x�A���r�5�P��c$#�f���	H�i�jk�]x��Y�"���O���n�^*�/�������iS�c�U e����"�*�>��?'H�!|�s�u~���q�OBGk�z�y��# ��S� �n������1PRs��	TD=_c�0��9Y���)?`�N���3Au�N&�Ip��ˏ��V���
w1�=��$�T��o��Tŝ;�l�>��<Yv&G��Cv�b����p)�I4�v6�z�q��𚅻�1��.X>?���7�?���l��M��zR�����<���Zҵkm�Ӆ��<>-q ʄ\Y�~�7���,�3����ab{�4���g�]ۭ?&�c7s�˕�a��]�.�3Bw�wͬH��������
ž/]����~}��B�	��6r�����6�/i��O|��mH�u^omS�����@N�ֿO����d���r\M��v��k�˗�V�0z�ȱH"h-W�o�_ɜL��'e5��� ǅ�F�̕$�x9�t�}�$Ef�t��i�9���9N��&,e�N�e���bӂa�y�(���	UCA{�rҠy/g���l9�`ڪuB�l$b"Dl�ᷜ<wt���*��P]l�ʹ]�Lj(eރ3v�?h[��5�%�	b�X�O��#4��Јݾ{M�Q�XFX�1nw��j)��k'D���\ x�N���ae�"|�D�Wt#*b⨲��_�>�"K��:��nJҺ�u�G���]x�Ba$U�����L@������������,JϗPB��X��P�]�B B��A��t;CeL>�A�^ob��ҖQ9F<��.{&ċ�,Ae�����Ҏ��^BڜGk��lӢ97���X���ϛZ3*sv��R�k_����V$��d��,��uh��z�-�R�p7��<�Yu)6ǰ�s��as7�X�rZ˔]�C��U���DA� `�(�`Qom��	vO�R� R{-GQ��p5��^ik�p��sAb6�3|�Z��M��VZ}� 
�q�g�r���2{�2��2u~UPe���Tʉ�kDsYl\����`�>jN�5c�r`�Ó�h*P�n�űq��]?<i��D�\������+�3���@@��Sk�)��>������\:�S���".���=�JM��[h�hwothM�s�,9oK$^��Y9gD��br���B8�k:ы������X�3���T;'�#Z��,R��0�l��7�0��f"	Jɾf����&��9���l;}�t�:��H�V�Ex�4�S`"/
��ݷa���؜�Rm{M��k�?Ԇ��1T��/�Q?����[R7.��G�`�P��i�/���@Q�CږM���Y�	g	:��^r�{\K%���d1�	�m�BAL7�bp�	�Aƅ�^�%,�+����x)�=OX���xS!��~��x�آ�|Ty�uh����Ψ��Q�"��m�[hX+�q����y����L�Cۏ	�>wnD�oGE|v�񼜊�-�1��Pu3�0�rB���3�q$5b��7�%1W��+���k�7r����?qO2(��r����\7(�u�eb<�ds�Ǐ׃�0W�3�(¶��5z��F@&���t[����*!�[�=S���ή�� ��-q�+��ܡk_�Q���{��)x�g6���ZD۪\&��(x���B	l��hLy�V
E����	6�P׎~������j�^;�[�T��:��ɬWў�%ӫ#�m�v�y81w��,M�l��|���0�4���䋟�C@��ۙB���@���*_��
&����[n����dja.,�!��,Q�N����$�넒�Y��h�|7�NTƍy���k��&�����$��$�	6��v��--{�(!�l�#���*���z�z��w����Б�)D'���	}$u7�;i�b>�>`W��/[i�P9���=n��u(9P�
��<���y^��@�2Si`o�'��a}�u�m�������X�)D��J�^��p�~��u�X5����E��wXm,����n�(�7b ��z��~j	�Z@�>�|5����ts�r}ܝbw������]�l�
��Hx�0���W�;FEp�aV5�{fhM�.(�,�1�'Y�L���n-��0��Rx�(e�=YfDf21�T�y���o�L�M�Vk�	;X�<¬��L<w�G#�C��I��)� �U� �� :�W[M������e`Û�Se7�78��B1S�fwtd�/ؘlz�5�+<�jc��HMvPbJ�ҕ!��� 3u�5%�PJd��	aQD�dM�� Y�u '��t��%4mWc������G����͆s�
 �eYX���FI�D.8��Ya�����K�����`آ��"Ngs̶�tC=�?�2-��(� �+�=���2�g �2�� > l�@u�ܿ8��Qв�M�A�
}s�k�U��?��'��m�Ck1J��I�/��Y.��|�!o�pyW`"B��M��"�كyU����b
M�X_���T�у�6���$]JU���,���r�Q,Ќ���5����4O.�䨳J#�O��ӷ����km��)�q�Mˡ\�	�_��SҜ��v�:�X�!����(^��엏8!���O߄b;�A�&l7&I�d-�[`�<Z��¿w��<�8��s�,��:�d��w*���|c5�	d�e��OL�]�S<Y���m8>Pb	�)'�U��{�|��%U��}Ԇyn&ɰ��8��Y��]c�*�����g'ː��7�l����H��n/K�ҹ����y��K�+����m���؇��JW�*��a������h�2Rzڃ)[_��͖-HiDᧆri-�����XD��l-ܤr�Y�ƈ}�Y�r��l��34)µ|'Yͷ�J	
��>����4kL��H%]��t��M��r�E5L[�M?J�������e�,��[$]��������k�mCn������<h���w�#�
T��5,@�<B9� ��^ٻ���O��ݽПbb:�ph�*(��5��uv�L����-�r!�q�Ǆ=�����wq6��@ϭ�ؿ,@y ��@��1��e�b�@� n�II��u�;�á;��2l�P�#���e)���ٵs<4b��Y�ڔ��X�If��ǄX�=��Na��p��w�Q�[EEx���{��rk�ӎd� ��w���j�	b�dMthv��(@O`8��J��e�z&$���溜�A��eS��`�p�n�rv�|p��dJH�іI.\!��U��B�����=�X���0��[|��������?���Y��l/�b����L���j+�|r&�<�6~�f��,4�q����"�,W
J�_%v�oT���Ld3���7�A��b���d��?�U�$2nc��c�ԣ�G��\�{�Y�d�F�q�Y��9��]#b�q��9 �!l��%�x~҃Vl����h8�B���V�T�u7S/�6z��8��tn��e�H3KX�4�G�����H��UY�w��+�d��0�"���]? <���^�)�?�:կr��1����ػ����Üﬔ�?:)B�UQ�ƕ��d������i,�b��ܲ-�~���@���J�9�x乓Ѷ@�N��ܖ�֡�{PQk��� ���H����e��75�#&��a���1���m� �������mE�řF^�1����U���z�0�Q(8���/��,��h��'�	�Ggs-�ޜ��"��se��2����v��;���*{��x�;�h�5���  ug͕v�R� `ϸ�7��sW_�_@��~�V�g������g]��W�Ѭ��?5�L?��$^t�K
���2In����:�Ws_<H�F���}t}:?��1��:$�0uS*v�Q� )�4>[�.4�O�%�N@�.�+7��W)����[����w݊5�2��F���OY7�V��wp�����>�!c��H��N-*;����å%Uu����!7u������e�=W�3̈́3�/�ȑ�XU���ݦy��/��[��-/*���+�ġ�����I�`�O�/���Du�lg�����4�R�-G�zz�OaB]}����֤��P~��F�����'�7۫�)6q79ol�.��� l�6�7��g�S�ɵq��Nr|�MA��)�Z޶�/�~x������ȯ�ݩ�+���#��u��N��pOU{���(�m0f�B��4^ߩ�QH��X�?N��!^�z�͘`ql�y�b4�R�F�����{��R�Oz��-o��~IV�c���ھ�.��S�\vhCe1�u���۴	���Z�$AR�������x�%Ӆ�#�mno�E�R47�j��,���G5�X����[l�R[Q?zMf9��~��/�c.pk�����N~�x�S񊶹I�liZq�����)�E(�2%������]�	+���,ܓ��%�d̨ͳϫb�Ȳ�g%Xni�L�KXJi����T�E[ڌ�Kp��տ;��4<��7����}d����J�&��/NJt<R�7�G�PfV�/�	n����3 �T�I��Q���2P�^��녲e��3�=k����:�P0� r&&T��s<Z��*c��$K��^+�ӱ� .X���?Cc|�I�`�v�w�D�R�'�b�!��t��\�CP��0A���K@��
O�} �E���c���S��	a�����|-?.3H�F�4~�je!Dԓq6�=P"�n�tM1��
9����T�a���u���Eէ]�q�@^��SO��AhQo���+[�x����c�7�fK�Z���z�|9S�0,-�}��{�+��}�U�H9��'�%���8A�௘u���E�|-Db���`��[uA�h��X�Ͷ�v���3i��~�p���<	�ud�?>���s��K�p)-�s)8�UϺ�f_BCT�g�/�[���eM�5y+{l��k�TnIC���VW��8LX�_ԊP;!�X���"�hz������\���Xԓ��;� 0DF�$���qJb�H3X3���g�vo��lʴ6x����q������?Uy�gjp��NAg�zebT.�[��^c�R5s��$�zږ��ؠ������$��#�v�й�����""m�NF2��!H�Ip����mi/�&T�3b,��IM`}�fGF1q� !z�̏���2�E��*�A�aX��7�#���,IٕN����M�"���I��\��v�>j���O�0g	1��ϙ�/�r�`t4K��&��`$��z6%���W�� Lm>v-�ʙ-�/�U�.�kqh���O������N�)���rH�]��$&1W$�b�ړ�'Z�<5�/7���Qz�xK�^pO�9@��=�1�>9��@P֠��nBY��K�=�o����}��,`fP���M�/M:�4̽l�mŊT>���N���\�ЖLG��E��&ի[��&�Ľ�'pBM����R���_���35E�Ww��GƸ�$��F�A���T�۞�Ż�C�ǺҌ!���{|��+��(����y�B�GoRŦ�6i�-Ч->R������Z3�)~)��2CHy�ud����t���E'G���bKΜ��L��Hlє���� BG�+P6<���2�>����H���&h~�<ɥ=�O���;�Ŕ�Q)X���&��^pG����Ė�z�#������Mcr�L6F_�Q�}-�}��8w6��.��7ց�QX�EM��C�F���p�,g	m���s�yv5v̷�ua#�X�Me�uI[��hR�R�9y�j�h�s�4S�Q|sZ�xVi�
���(`�����k����݀�9|�J���k�CF��
�.[�Nl��Ոoe�3ԥ��y��b���E�$ʡ�8QG�j�s�g��+�����^f����fC!���}ؽ����SHY�U<8yk�d^�%�5��,7���6�<d��>�4(n�x-�a�������6�O��/*]h&�M�� 墭Z0ș�Nn"��	C'qwI��{�l���[�K�Ti b���q��,0�����
����ɥ����
���b�Ӑ7�Y��$�K`��(�")��-������m&-��E@t�u�*���CV��Z&��g(e������U���И?�P���3�ɟ9K:k�h�:�z� N�y���#���=e�r��}�="��T	)B�F�dE��~o�*$�g��*�솱��j����l�,"|W��(R{��H�`*��s���8*�Ʀ\��&3�<�P�Fzg~QkUPr6���67JW�s� � ;����!�Yeי�B���ث����M���E��2�҇����Z�
�&q�"-�'�=_Y+���*
�����C��sv���R9"^�֊��ܐ�٦���V�"�f�4��Pj�f��*w�C�Z�uf�C8=�����Gt�Ю�
�$�ea� g3�%��q���t�>�-OQ'����� �t�t�WD|��_��ǟX���8M�2t��lYh��I���4�4�(���c��VA��I�*TB��ͱ��{B���ݎl�(DWz,y��޵���E��$��t�_�����G��N������K�!q��Q�dY4�z����%;�
�L=�:*�i�o�R�Ti/�#�w*RD�:}汥F2ODZ�ʙE覍�-��E���$��a�$SI&�ke͞���ÿ���_!���:s����ŮD���g~�z�l�n�8��G�:�^��`cD��I� v��<w�f�Aɰ9�m���"pdRg�����M�E&&g������)!�a�9��͑�%�(�/�=�*��/	(-�4�̊e��h{!e����v��)<U�\ucO:�vg+�폴�!Z��k~�������,����Z���2ͫ���o^C���7g�4��\�����y�E���b.G���.��v�����&��6Ze�-9�s�1�T�"��:��(����Gf��f
گ���gjt[��P\.�&��x�*'='�gR'90&�	*������oһ��Mδ���0'uMAl�?�*M��%�8b�n�w��{B�����M4��J\�CN��{/���!)^^�Cm�`��93�
�p��N�⾖�+O�����&|��`h��\�kJ�r�خkrG� ��
?�츍P'(Q0�{+5�[3�iو"���1˔�g%������"r@��Ê�u&T.�����s<���)�Wy��K+�d����H��@
�j�;H������8 �����-���Z9�%'��
^����^N[���A��x���ѽ9�M����,����2F�K��7x�W�C�� #K8� �h�rm��b �Qr���:�?�77�NG���?����B�`�Fb���BEdz�����A��O���������{B+@�zX���*'o�/��
RI���[/�A��h�(iQ�i'5lػ>	�0��^�Ζ`�J��{�Vmbymt�;]̧��?%������L?��%u���JG���S�ܯ!.�����#��&Q�����g�gb���|ͅw�����Q|��(����-\@�C���u�R �)��'N8Ƭ���`��{�	t-z�eֲ�{�͇o��Ѓ����Jm�
;#B�H>��f�[M�[� (1ؐ,��%�<���k���n&-z4x6׍?$(ꌻ��]�O�/m�v{K|UC^�����v� �iN*�ǣc�ק�^���7 ��������9R̈�]q�~��>�
S||�y�xqqB~}�qM� L�V�Y�іmG���6�����a�x
�6�,�k�0����^��,)�@t���C�V��~T��@O��N��*@�Vq}��i�#@܃�p�4o�׆1�2��}�ё<�h�H�|��&�Kw%�u��C3MyΪ�DUC����w�kn��zu�����x��s�&�����Iu����y��<U'Ky��˰(X�P!t_�<b���s��
�μS �+�N}2�[TI#�{Zj�x#�'n��!���
�HJ*�P��ˎ�!�� TMS"�'���o!��Z����.x��������A���c�V9Y�W���@1C��7tź3��������D�U}&��[m����P�՟�;[z�}�ѭۖ�w�`~Ϸ$�E\E�X����� Yb���.Τ���x���p7E����>u�@��� �bS;�@ԏ��kw;)"�,��fn+M-��yw�R�)�jhဥz+~r?���s&_�%dg�d�.B�j�뾗���&���^�a� ��OwT܈*��\�����<�+�nw�Q��(6��f�y��vd�p*6]���ݕk/N��9���"�u��k�'C#�:L�fF*פ`I��"x1�r����2���{~�]�y�@>1�%z^!�{�'�_�*2�|UI��ư��3^�="����q��)���lBK���m�/��8��U�}�ymjX�5���D(��Pm�C"+FbQ7�Mt]�!�W	����4�@�H�L����!�u�D����mw��3��%^�����w����My���(��q4�؃��d�z�����@�Na�!��É��g ǟ�,�u/�\^q�p�ڣ�d��zs5G؁�����˭a�KSd,�,9ݼ�U�?���i�E�(�H�YЋAs
�X9�D}�
�a��+!s¦|$�D_:Z*<>��L�,��n��$8��8�iu���%��Gn�TG{��[�7K.7A���|Ϯ=�3���Q����_�&�pq�G8xR����x��w]9?��8(�'���7~G��zk�OD�	����2�]m�4Έ\�?8�ȆG�wL�gv����S�
��7��yr���N��[�cuC>�H����(�(]����ǂ�OI��F�q�!Ai������K�D?��'	��� �k��ri\�"��z2q�,6+�X���ʑ�h��u��=�pW�ԗ�1��;�\*���V�������!�|w&���8S�a��=��a�L�m��j�C�!5~��ճ�[��Ѧט�����,���Ȏ�r��va�c�٠�V��W�(A|7�2�/b���-��L��>>�5�(��O<�A�z\�S����b��g�XGZ� ��=�T�W��{��^�|3]:صg��܀u�է�7wI��8kU��m�������@ՋN��b��5��@���hkk	�ix�dt>�(�2� o����j;,B,	o	R8��ѡ���ʸM�_�N[��{#Z*��VB,�oʣ1�wF���U���w�g!q�
U����M,T{P�x �^S弛� ���y�XD�_��Q�W�Md6Q�ބ��sE�WQE$�9�>�xD� ��"n$��;	�F�����|�����2�2��$����_T�x����|E�"��$�3�Ѹ1��_Q�I��˿�����I�gӋ�G@A��|CR��Ie���;������{;�M��}���N)V�2���Wpj9���}gr�-��c՚i41EOY��t�p9M� z����[e���hq�7�V"$��hą(O�@ol%�"O���L�-�hv.����"aK''� ��,�I�y(�TaL>~5�4{�7��|"N5R�V��ꓺ8���^�����%��g��r��[�G�v&��Է���\�n�>��GξDH_,�/0�W8�� 3U��b���0�� �Ў�������={G贻�!"A0)�9��\���*��E�� �V���w̅GoNe�x$\��(�ɘ�Y45���s��"O����|x��q�g���f^�n����]�۫%;n͌�{I�z{9ϧ�x��y�9�H�iZ\�I�hDcO���[�!�9��T�����UM��1�7NY��� �ٜs|�������q�9xN��R���JɭD�M�er�I:��./!d�!�ѓ���EO%t�	H]dD�̟6� ^Z⪊.|ơ�Ϛ q
͖�j��s�6�U������6�nKA��/��1O+�Y5�3��Z�Li��?��M�iM�ڹ��kȔ�}gM�u%�S�ay:Ѣ!A(Ω��2%vg��f>�'�dn�ĕ2P����_��S�b�X�m8w�}�F���{�;��x�ޒIX"n���3w#�ךP,�	�����	��N)	�e�3|���?�%��
�.�Cw"7ov1MW�)�h�Iō�g�fQ��[��;YVȁ��*}�I��e]:�%�a���q���ݦDM� �1�ifq����i��f��gܻp��6�x����/Q,9H����O&jM��j7��WD��^a/-b��MQ0)�w����Sn�H��!xHR߱��<�����e�Wm,��3&�	�&���~�������h��K����l����-
�k�$���rYi3�R��B4��؇�&�%���F<c����	�`�%7�$~W�`�����MH�>��)�(ѥr�6�F���bsy�Q�Y��z3?6wO�qR5_ *7˲j��|���^��Y"�ֿ�\l*+���~hŪ�f���E���m�	�P�o����?��+�s.��s�y�t�{��Y>��;us�:���	7Ӊ:�o w�w�z�D
ב��e�<¡ u�FOb{#�Zֵ^�����QE@�G2�d�<> \K��ʤ�� �U:f;���)9X;z����R�����!P�*���T���K�y��~��,J���86/4�i{���1���_�g�>�^[��N�ãl���=AS�p�K���/���c�mq�q�^��+�a9,Y�[3�-����w�;�H�	�]�ƧJy���7vJr��(^R��q�e��v�����u��7�|s�o�%��QhA����j��\XةЪ3�2n�`�+F�K|!�˝�G�@�G�Ο6�qw��4fl?��ޜ�.�����*���PoҎ�i�'3Wid�S8��㖝��</�L+�`�y�/d�j0U�X`8��+$�*籠�P�	u�;��&���F��q�a���yq��F�j�Qw��'�	�Ka� �B�A7k�0,��|t���E��n̂�dy�J�=��>3�s:�n���?E ��R뾣Q�=����jj���,@T"�0��/���2���}�j�es�c��:��-�U���T�����$�r<���I���"��h?��p$D��*�7�����o�	��M�w�\{��M�1�c6������t���y�~qM#�`�CG�/i����ڛ��7jL�jvҚMzLn�Ƭ]��z!XrtΆ/�gGO��}��t(]�v����͉ �%8���j�m���	���P������=$DM���O��0L*��Kf%��v+�g�ͯ���8A��c�����p�Ϟ���,��kӍ;lM�4�)��
CR3y�YP�hre�e��H����3�\�K|����绲q\�.��im^Xմ�0��rV9<�]CT@����eÎ����ꁟJ���nѬ��8�k�*A�2H�j�~骒:bo��yẹ.��t7Ay�O�J�����@Cy��H�,��O>}��0cN�M�!�g����b.!զ�x{����&��+M��]�98`T��	]Ҵk��"�}	:�S��Kb�"i[����0B�q�� m/�r�B���[�֥�N<�]����g�w]"E���n�/y��9���`�8�'�;��$ψ&�no7_��&��צ�?���2�T�߂dS�j�$\ڔ��\x�����M���L�D�	�
�W���p�ڋ{����y�����D�#�r��C����<Hr]��";���ʹ�E���SG�$�����2�$�62���=�
�����[�� '��go��M`�itV��c��{�e6�f���p1�#U~�H�(�>K��;�^z$H��,����÷�^����@'
��ڷ�-_��&G���>R��\������Y��u?L�E�R��ރ$�J@e���F�l��f����5 Tem�$Gcr����al�58oހC �J�<��S����"�u�{p٦� �CızE-�x�}e�P+�yߍ�&~�����=�m�97��y# ��Ó���E4~x��Gt�Q���Yd�LD�:&؍9 l�4��!�����T���~LoW %:�ug@��|�+��_:_k��hd�,	Z��ci*�I����'W4�����gl^oQ�� ��l4��Io��='��	�n��/�N�/YR�x���sP�M�	��!� n�u��A�<!���yڮ�H)g��1�2�I�����[�dbw%;���}��w����Ⱦ�:�q�O��X�<IŠp�YA9�B(	�9�������q ���툧�oA�5���:�^�;�~YuyFJ�?_�.�N���$�(3 *�W����F8̐��rx%0���@r>c ��jF�p�<٠Y�o����?#�պ�F���K�(��;F�ĺ.�%�Z�Sg���<V�Z�4M�L�����]Q�ӼM������RS=�I��wQ���Iѷ�c5���U�Q�0�N�wwn�yi�	���P�G����1r_�6ם5��~��Fj1ޘ��h�Asj����κ���1��*�����p�A
b�%�ϋ̽"�0�@���Q�����3�#1EE�e��J�?7��E�Ϗ���*n�P�	�خ/����.-�|P_F w�B�Eh (,GZ��U�nu�n| ��'(��[K�Y��N�dd^�5��g�`|�^�������%H�-�I���<�B�,�=y�7�ߊ+��GE�:����}B��P�Q!R��-YB#Ӛ=�[���^9��W�/��m��������'�}��+�����b���# �:�������b�۟V{�{óW��v�`�X���1	��I�Կ�M��g��@os-)\�?��k�����&�d���r,�0�f����6O�]�g4��#?�>Œ[-�2�Y� cl���Ռ�'��;�����n��f�k|1�j�����(�	6�W��J\�QQn��ё�u���2y!T�'�X���5'e���!�5^~+�TQ2��1r�߲��Tf���H�����[���C�1�T���>}�d;b��gO6��� b�`�9G�Ѱ.��وS�y�x�\��l|�-V��[I���
�z����ŏ@��FO��a�(v
/ڔ�4�q��g�'���1�@[�a	?��y��e�w�!P��"=]��,��݂�Qo�L��֚��ր��֞�1D=	�#��4���!+!2L7T�Uy��ە��Vn5���}_�ײ}���`3 �SgJ�s�^�a�g���^;��Ĳ&SzV8��h�I�$Fi^���8 ��C_�� ��X:���"'�#Kr�Z��r4�Xl�_M�~����4�ܧ���^Aql��$��ٙ{��mZ��vID��l-L�0�x6uՇ�%@+��S��J�*ɔ]$hHOG��fNyݓЉa-�W���-��UA�*F�O��y稤����g#L���S�~��'{Cr�@h����Ϸ-H�U���v�/ܦ^�2�J��so������a�/��MM��
�O#,��E�����蟳��\R�L�*���2��a1�(B�.btT�x�:OcN�3c>k��n������/��śAR]��_�����<P�貀�op�P�>Dᾎ9Q���~c�������+B4s���}��ԑ4I�$�\�|�h ZN���>��G#�\��}:�\cy���Ǎd3m�>�tx���r̷��AP�$�%�b��-y�����/�e���^>�Q���Rc��O����~��IV���#wǞ�i]�6`+\癪,��kM�b���g=ue�id4O�{C���G���=s�E<;G5��7��e��w�z;�Cm�;p&�]~5�7�>�H�и���I�m�b������Ǚ��嶟���Z����]���1�n;�����=���� 4�Z.05y��U���+���_&�W�W�gKn��K���ѽ�p���)6�8���$/�Xvv.�$����sj��:�(���z�GC���6K</��`+��$��[�`;�I�9k(G��!���ت~�aX���|9�1�� 6	�@i��܃Y7��Kc�2z򥪓�{Q���tv���e���N���4�rޏ*�����R��� �/*^�ޠ,E�oJq��^�־����oU�D��6���y��$ʵe�~}���-��A�кҌ���<%�,�&�4��(U�d�0��B������Y�Dd�x�C���D%��w��N��NCT��XŤ֠2G.��� ���֬�.�4�-S]�M���X)/a���}9�|���e`nQO!=�r:i� ��ݺom;������_v��ۣ��8�$�Z�6�'��
_�لkT9�Z�Jೞ��1��>b8���(�\q�{�$�B�`������(����Bʠ�{�^%�`NaUe�~N~�GCw�cư�v]ƒ�7{� �D(&�PG:��X"��n�������J[\gaT{�Ƶ��ٜ_m�4s�߂^�����+QgP�:��p��̹���+V�A��ߧ�?��Xǜ��)���veQmJ��)vqw�+��['��\���?�TuD���^
I*IWqS����rD]��-�. #a0&���e�sɵ�1�����[�;�P�������@5y=M�
h2"��|�������8�m.�2����V��B��F����!��̙@݁`w����Me��A���s}tF��tRmu鐛X�vo$�S�I�'�9y!w~J��5�I�����4�=�W��#�?�D��i�p&���y��M7y���Ɉ(E�����{)�����\�D"b2��u�suV���*(�݋ݑԵ�nI�D{�<��"��T��h`b�#_����J{�400�3�~]�n�9��S�yP��!���L�9'���M��ph�ʃ�����w␟�R��a�窒��ԍ~����Z*Ĳ������|�Y:��cDm���?=D�\�����o]�����	����{o�OӝE���V�l���G4irh_?�*%���Y��f�ׅQP�!HU#���]ek��3*
��~�6�,	��t��޸*mOr:���:�
���AV�u�>E��Q�?�?��_�?�#�kq7�7�3Fy8�D6r-�G��|L�9����J�;C^�f<z"	v6��������޽Wx����KO�Z!Z-؆�55'`����/g�	���w҈+>3�}��ɒ��	8��/�����}�0����=1��ނz�S�;��#�q�{����=�;�R��z���wk[W�����{,�����d���E�P���Ū��}w�Q��Z0��AFޮFܢ*p=���[���C��*v��N��Ҥ$j��E�_o�/�P�wj�0U�dd,��?4O��_�T%Ŭ�J��V�uf��tD�ҏ�����d���߲y��2�H�M=��ק+�~lkelT�R����vK�p�۽�TPX���%��K���j��Xf\�	AK��f��@H���� �����WӠ*�e�|���`@�b���k���}�nm�N�Ү��(w�X_��?�'klWQC?��/O���@Xb��ހ�i�>�C�:@�$0H��n�����E&mly�P��V^A���?S6-���j(`H20L�nO�$��!a�����\�K L�_����r/8��H-%c�*������i�� �'�}���jL�
���t&[[��s���G���染
˾�I�d�b�'��<�s=^l�"<݊�����Sw�K�I�J���TigoXU�'�7���Իs�28��$��]r��H����!x0x��#�q�T�@1z*�q5�}����ꝍ�����Ŕ�=Ω�%��~��=��O�7U�MeE���%ڄ�3��G��9z7y�^Zw�����n���P�x~��W�s�?l��a�~�L��1D���O���N���	���$�|pgy�$i�$x�ʬF�է�nPuj�}:������Z�Zz��ZejIvY2~I)�/�P�{��`)�ƑE��>��M��+p8�0z��y�w��;�ňT�j��9-��/,�f b�1C@e�. �iH
��Q��uK�����HT0x��Q�@��g��-}ސ��޸�f~ u,�jQ嗁l�����ڂ�;��R�����KOQ?�!���jw�ۏ$��fl�Ȫ�%c��g�{��t��CxK�Thl��T
ip�=�ĥ�a������h�eFq"�RlH2p9let܂�k78X��ؖ��#�D�����F������7�����F�~�6�����,�z�~�m"7�B��AK/�WL��U?Ocj�45�j���룓
h?/qv����f�SD��L�β���
Ȉ�g/Ux� {���8պ4�H(���I�&0B{5ʽcۍ�TX [���#A��-luD��J/uЄB�[���C����-"T�?`�"����{���eE����dw�Ɔn�P��@��
��N����K�@�b�gHJsƁg��xg��+f oO��K�"��A�ZtB%X�W�	��f㮅f�]��7f�@�{YM
��rt�m�M�0��
���h���-0��3��3�����t�'[l�����x���A��&�F@3a�SJ2#c�V?����YTr�X̒�9�<~J�[�X�U��Z{�wl�4��ɇ}@�T��ޑuԔ�wk�����R�ؔt�^��./w׎�ELrE�i�0�i4�+��	$�+1]����.������ԇ_-+���41 ��Q�@�&@�#o�B{ }�3k{2��
G��)��/O����N"�/o{Q�{��$�e��x��Bh�2)�$El��_E^�/\�VȽ�J� ��h����h@�I!��N�������hy�N�G�6T8�AYo�_�L&���PҀd�M�;1����!)Xâ�^�T�&s���í5�4�T��kOO��ON�}�2@꺿9�s�3��k�`�񾬖8T�6٬���%K�F4�t��N� a��O\��ƣk����x�����u������y_���Ҵ�DR�s��e� �E���o�M�s�nCN�E.��l*�q���X���a�(���Y����=��[��_���sv�=�O���˨Z��h�8��/<�@,_��[�J�Wm��0Z��.���ς��yd���?���834�n����ɪ��)����<-���`�h�,����h�M�ʃ�zna��p��@7���Ÿ�4�d�^��Kë}�����gb������N�*QM0��\�C���VeU�6�.����B�I���a�v�r�^s��S�����&��]Wuȉo,�pR�\��
Xw�E "��
�魛S�6����X�{��1�ݻ�������B^��E��+��"�a����>x�[t������W��'����f~Pz��B~�y �!.����p+~�|X�e5�j>���1�²��br�)��5;����ņoI�,���QПc]vn<+��������	��{�L�1+����"�FE�|I̠��F�J!���x�n�s�OO
bN446ڰ�
��@��я'i�lѼ���N��Nzylnf4&�L�����Nr�
Q���y��7%�:}#� �!��`b�_<���v���҅�s}L2 �	K�z��d��?@��ٌ �9G g|I��y�"�b�X?s÷������|e��-�e��$!�%t��EX6��?
k���7А	��k��S��)���/6a�bWm�W�+�k{�B1��%9N�R���M�i�j��n���������:^���ǖ�S[�<K�cqO�\��V�4���IҞ��J�kfQ���⑚�O�f�Sv�Bd{�zZ�0���3CZ^�h�
��	X���{�=2���1Ͻ���z9b�fk((U^޵2e��P����������J��|i�߰H�q6K�.�6P�!�x�ޝ_�A�f��l��%�QD��w�������Z����36RNe�8K� p3%�żs:������#��w2`
3�̕D
��R�B.7�ֹ�vk�K���@l�z�tL�v�"�23xtx�+�];+���\�1������X���5�Y���"D2�0ܸ%7���ͰZ�<�0QNG�����MyO�|��m\�D�x'op���蔛0�6���	p�vY[��������:�@}�.Qdꮜ��~+��@��r��h<\S����Γ����ߒ�W�w9M�t5��w+DJw�2>�R�Tf�z����<�?f��#�/�*�^�l-U�=ߴ�Fg)O��ـ�<��c2�}�vkK�xX�����6�>��kpW7�}��{�]M�׼����գ#0�z�61����ToY�c=�I)%gmI&J.���00ylR7$�]�U�e�9���K�Q��#�-yN#MTn���T	�?R3>d:ҙ�.�\[ ��)�@f(�u��KY\����$����k����t��c ��sT|ɋCn��C=ÜɇZ���,��{�c���$��Q$-�l*� t��q��c��� �o9���ge�T�F'A�]_q���P�;[ޞX�IW�� S�hӀ�ҏ0���I��Kk>�S 1-�˲�Dm:9Wu�O^��h��0Y.lѻA%I�L���Pܱ��U���8���������0�!W����}vs�Z����J���B � u������p�*de,��4.����	�F|�o����ѵ̝���rݼ�7U�7X�I� �B�9m��؄¬5���k2��ʤ��]�?���k"���̋}P�9Iң}n�BjVտC粯T��&��Y�1�
��7�u��*��������RI����C�sw��Ql���~��E���E�&����A��7�٤Y����B.j�!j�C&ב�+�fA��aQb]�~�����R�w�^m�v���Y��{x���`}*��%��-y�?�2�~�"�)3����NۺwR��ֺ!��r�8�ul��S
c
O�6�ɫ�Q�7��`J��:�ȦGg����ĺ����cwu�|��OW�R|(�ls�@Loz��k����� jJj��v�@���o`��3�e�
��CQ�Hpշ��,kd� yy<7��47�a�:RA�k�;d��:+����خ0_ڌO�C�f�u�ņ��::T���ZX�lCLrC�֊S����R4�fo<�aA����F��q��ʽ�� Ae{Ϧ��B��]�H�nd��#��#�6�!��$3�a�>��w_��̋N˧��\@-*����Y7R�O6�Ѱ��O��C�8@r��2:���'���Q�e�؉�\�}��hs٫�pW�V�A��O����&g�����R���)й�5��~�ۨ�/�?�2�]���}�5=��������;���wL�+=�s��zF�ϩI����dl�ˈ�tP\tG/-^�H���x�Ƒ��n��1�/�:=#����=?elگI�v_�> tǶ�~���%Xó�زP��6�ߢ��<���#3�B���5nG��t�I��R�]���)p�&�ҾI������oy��T��)��M�`�?�a�}&�P�˖����~��r�g:�b,�����x��"��d����\U���_�zC
,�&�Kj���%y����L9��S������: H���9�y�7���-C���r�Ó�g������ w�ZO���>SqK�O����l�`���\�*����r�B.P����]�a�.�:"o0zԬ�AKw=���uR�H���X! �����������0V���"������l��R@pV��Г���ջd�˳B�o���e�m�hGGV�%_��<#LL���u1^Iw����m�	��74W)�o�0�B\}9~���"�d�y���U07�"z�=''��-�v������"\1@�7|�F^�?�1$b�b��(�9s:L�%��_��qi$�l�-��A���ir�g����C7�V����КG@7@�*�����8Fd~Y�r�J|z�����f���pƔ�Oc6��^����+Q<�-�m�M�O�A��@=d5�5�]-�N�����Y��l���� ��F�0�+��{��0r�U�)d47iu�ۡ�� ���@�F�/r�/ ����:Mb�SH�w~S�6�?�I ��Ǭ�������筰����\��R^GB�H���X5کg�^M��$�l�Z5~1�5��8i(��p�W��E���8S�'�3�.�hx�Q�.�+[�}>���l1\r��~������.�JW'�1���;ͯ�]Fd^���w�\1G:�'~K���2	����'݆%F��uހ=���Q][������\4&c��貅����ю�Ⱦ��������(m�k�;f�K����\Ld���8����Ȧ�2��Z��eʾ�Y�;I����\����Q���8���?]� h\�?���$�5��,[�'��DIܖ��h�+�a�$P�m?0���S�8O&���E�5J��k�i�R��K��� ���"���Ed�%ZO�׻�|07%�J)���:ibp�A{g�i�Y��pܡ�>hZ��!!/N�Ң���(�h��2����~��iN�+FQ�����Or_qW(�%�S����]\Va�[y����%?�.ҝ<�(n7%����m�	϶�X*�O�N�՛vKo�>�䫿�fp�~�N�m^T�1hZ}���[eN=̀$z��H2�7,�62h��eL��PGi����뉽~A��}v��?�-F��D���^s�)�-kc�����Y5ɼXK�Y:����c�0�Q�$��&��"5��cUz�Hv؅���"U��x#"
;�6#�[:Ը�K+�]���% �~�� u^�b�m�Lc�ƴ������j����R8���H����&����S��v�'}Ȓ�>|��X�<��l�ȹ6k�y�m�!��]6f��������S���Q!������tΖ�5��!��8WI��� 4�'ߍ%�{�9�6�_���6oi�;)8��]���f�QLHv�p�˼b%s�n����z�SB^�����Q;��aTlȣߨ�'��qo&(�-�c���R�7Jh.5�_�)ou�Z��j����9���!s:	��~�Mc���
"�@�أ��ƫ�����ճ#��f6�=o���״�'��n��=�=G��͂��wV+w�W}w]|�z��t�:�䄌):MQz_��mzNu����e��س�x(;��7}:2��e��������y����m�� &4ZG'���<H?$�΀���C7��r�1gI ���$�YH�w�4L��e2p��0%�g��,�u�,�Y�
[��+��:z�c��(�����i����>1ư�*|$z2��������](�
��" #Brƭ����!�tm����Rg�'��c���S�
������L\7��&}��<�} ���b�~L�:8�%
�^3���7y�qCq�D*�s�h&ե�˽�>�����ȸ�f��<
W��Z�x<����h'H-��;�v�')o	��ju�4R{Q�%�&��������9��f��C������������Q|�����#/��SB�Ll#5��7nv=���"/���;OJ�˙��A<t8aQ.��A��d�O*	]�	�ҹe�um��Un�l�e���]���{?����f���е���C�����<�f�1�s.�N��_���JA-��_f-1�%[$3������ӣ��Ǣ����h&����ۗ��5�.x-�|Ny�R�v�%��/J������_�+=a:��{H�<�`� �}SA������>��Z^�j
1�V�~o[�Q�l߸�<���/Sfg1��E��X|��ױ�޹JS���mNB���]u��;'��gOC����ino�B�0!7.���
��o (��ಮ�t�M	%��� F�4>&��(E�~YYY�m|CB��)MG�Ng(-�X� �b�RͶ���R��o�)�"M��ޫy�t��8�V X��=�����G.8��m���_w���^��]����n�_�.Ȗŋ���J��.��C��,�<�m��V�l�{;�*wHKg
{�󐞁�S+ l�y	�`���!�$������Q~L��5��Fԯ�>��Z�����@2~���D?�bDIU�# d��2E�t��I��]T_���=�|+����vTc�k�[xSN\�SxA$\��,_�:��vs-Z+�b�e�@�w��_Mn�fŞ��_%|W�_��A�UX�]���3��w+��o�t�0\j0i"f����O]�Ӫ08���~B�OϦS>��mG�`p1�]�a� �a~���p^`��54�g� jn���/9J�;~��<�=�����m�W{��C��DQ6�()	-$�p���<���>�H0	 GM*a�AM"���W���U��3����W�L��cx���5p
��3��D#���jl�i�#-���|9��Z:}>�K2�KDJذF�G��18�9N%XWB Sӡ1�u�û���]|�_��}�;��A�+��P�9��o��V ��]^��SgwL���pp,5�A�}#���)����tTa<�:و���~�@O���[Z�2��-1��@�(j��'�ׂ}�顴+�8��2�wL��{?�B��t�OVP�d�ڥQ��\/{3�!�M Ŝ@��إ�@�V��Vx����2*9w8��%���=>b�Ϡ20Fa��\β�v����4������n_Ha'���L���!?xtYR�P�B��eg��e��iCX{���7ɞ'w�i\� �bH�(nT�\��(�+Ң[a�P�g�+��D�Ȇ��?��/��ՠ�Ӧ�	��N��V������3&�x��l�1��Mg�^���.l�N�p�l��fF���f;M��E�.#\��)�{�m-��~����fk_of��/ DT{f4���,X�Ŭ������b���`��M(��o����
�������*mԒ\O�?�J�(��)H�e���Pe�ّ0o�>+4�Z�-�׾JKH��&��2v�9�Y��ȗQ�u���PIY�K��gF������5�[uO��'���d��ÅM,,�J�̥<�W�������\�>5�������<�P���/�7C㤏�ݑ2��~9Ǜ��l�z�7-i���0�B^�b>��}ц����Y�H�m0��Tu�X���s���<���Δ���׏��[�����5�NX�v�Լ�lW�Xȍ�mp�	K���,���C#�CL�IMʖ�(�(��zV��Mwd��n�S�]�Wu��&�����ˢA�Տ����:=�i=	�<��Vc�S܊S7����!Ű���i�\�O������Y��z�	�{YX��m��j�����@M�Q{�,���v���L�/l��G�Q�?m�
�.��i픅�L�$��	On�&�/,LW[`
��ϤMt��F�K�/��x/�k.����Br�ǭ��?���ױl��y{�f�zI3S���>L"&���'Ve�!���M{IϹ�N����c����݈�EC?�T��*B7Jtv���6�گ��1����h�m�"#��*ГUI�c8,��}������t��;����k���J;J�'Q����B�E2�a����އ�Cln��?�9�`�5��$� ~7���F	*2�RJe�n>S�K�:�#h_5 �?�,1n����'�?�F�\جMAq��y�񘕽�]2���\W芰��τ�ډꑐ���G�
<(���"t��
?�F�!%��[��_Wy���d�Q8�����w�e�3��П�_z�y�V❉֧��N2Wz,;Zt!�/*s��$=��R�[A|p��n(o��P��0��vdF�Y�e�v�֛R�`�.�= O�("�A��ܭ�/*\�P�)��O��{W��Q��_qx^S��W�>�ޔ4��x�.F�/`(\����*e���Ǫ��ZKqt&��+(�n�9˭Q�m�9��tkuآ�"֩Q~K���~�)_r������W�
ݯ���ƿY�p/��1qv�J�Z�_��׳�u�5�	�ބMI�ݛ��[\�l٭���1�7b��#컍�������-0�ىf�h]d�sU��6�mDVM�\�<ಽ��6�=`S�J��Ȓ�������~B�ls\`���Ԃ��D'�q�ύz-��v�>��T�X>�|��Bv��Cڕ0�4&`��_B���c�Ӡ�]Mz�F���ι�Xo/��;��o�M��$:�W�B�W�@ !2ּ��'�{g��z��1�?W�́+I:�kRepG�B7?R��Ʒ�L���E9�Ii^ �s��Ng6�U�G�m��Nz��;X�tѓ�i)W?�{���c2j��>�L���th�N���C��mĎ0@=�n�kxd�2���l4B*�[���l��$����^���鱒AȻ�:"8ڋ��ؙ��Ǧ�Ei�x3�=�{���|_IB|*X�Q��X�`i�'�_$����MNޚ�	z����+��[�O�I�n%���e�I�S�Ǝ8Ju:�O�<6'CFh�S��D�\���;8+S��A�Ҽo��f�����`V
�_����44QY!�>9<՛����BD�.EEd���������˙�s�2:��^��߽p��u�x臭x#\@��z� `�(B��A/}.@�y3��n^�v`�r�����-���c}Ct��3�f&��0
>q6�������g�i������(����>��-���M�\�x1�q�x�q�6F���Cr����i�0��%<M҅Ģhr��D�ꝇBh���s?j*�ߡ��i�{z��XLuN�_]���3�ԯ��_e�T�ӎ����Z��<�vq?k�ո� �q�۹o���d+佌��UH���U��H��kӘ����kLLj��R���A��� �h~���H��iBz ���uV��fƝcvM
�<��* B{[�Jk�pq?l2��U8��HJ� 
l?���7�ZD�&��%V�hO���Q�/��B�0�S�vF���� �IA�����P��Y<��3��/q���iKu}�p�P1�w��f�K%GG�ޮ���N��yθ7���Q��ߔ��tl��y1%��#Mޓ
�4�r�
�g4�F�,�oQ��fΩ���&�ٓRM��y�he�	�kt?y�8���$Q��!=a[6�)O�\}�7�z�[��g��@FV����\�	��\Z_y]��Um[NUs��V��v�&��Cva�W)"���W�� ��j��&���:�1���������=]
6�%��;2�L�>0��gc�*x�z_T?a�rN�WC��_kD��2�7`���x:�OZ��zE��L·.#\-+����$0��Y����7/�)!k~i&3��erJ/|#�Ȝ�S��՝߷��!Ms,&�-ˆ�޸���?$Ԏ��3%�X�zX���O���~�:S��n=��|&��6�eb��[�8�l��&�1�fyE�5�2�&,h�ǡ������;�ߒ~�__� �+�&ã��Ա.V-З�?�T3�`,�<.�C�g�n����+����9m�*�� �X��g�!YJ�o��<a?+&��V��v�H����݊��/e\�VNiB�*�����3><�R`�r���1Β�)�Bz����O־����f�}|���*;�>)���3���9<t�9�0��BK��[���|���u�a��W���톍-BW�mp��UsE�T*N�m:��m�h���K���(�UɮQ�&��b'V��]H(��:�P�W�9��Xd"���w�T�-���N��H��!���I�o��Mt?p�+,�3�}$持iM�]��Ҷ��f�D����V��GG��\��)�X�Nq��>���~.p"$�r$J�(��U��_���X����\}�R;_�~�lZ� r&1���8%Ρ7J2����b����x�г�}��x+�4O�	�3aС�DA�i,�����]���բet�z�=*~�l���Ťz�A3�x�/{�Ѽs��h<�Dg�@�W4�IC���Fϐ�9�w_0�{�8Ay~-�:�
ν�ĩϚ����C&�d��ý��Xf!B1Hց~�e�CX)��?����j��3��X��W��o�4m	�1�1G��ڔ$��֩{��,�g�������m4�aW�q)��p�b�0YK�:N��k�����)lu=;��̷e�-���!��$ � ��
e��;�)��y��UᴲPi�J�	��%,���4�~�����bX�$:.�ʽ]7[�	��V�9祇(r�ϑ��7r��6[v+�w�	�����< \f�����Z1�ʠ/c�"��;,9|T��N!���	O�77���Ǳ�;i"n��b� �(<amY�*F1:�>��%"֧�%�;�p!���?47��>2* ��*!+�j�v�`��|#�֎D/�!���Pۦ�[�~У�	V7c��w>�J�S[��1�w�9�6��mGl�C�]���#�D�Hy�9�_K���Ny�\dy���ۻg3�x�MF�P����.�	X���{kAiu�����?��9O]�g����v�;�7D�J��/K�1�;��3��/��y	�
3--?�z�?���+�DZ#$�?�ML;���xDA�l#YYS�z'sbp�cg�*УJ��.?���~�_�>�:��#r���/��_�ԁQ�cY�l-kx�i\�;��УRm��o��0l��h�'��e
��HR����,��XZ�̌�6�Z��ȇ!gC\�j��2�`!A�-�*&`���ԽGE���Kc��sU�A˖��J'�9���~	���F�Ѯu$���0r�$C=��#�nxa�צdlYE�������V� +� ���!T����S	$�5x�jPA�ط�z-���<�Y�Ӣ~s��H�❂�m��*T'l����� ���-?��E-\u���(5a�"3�' �
Õ��RY�l) 5x8���MoZbL�I(˕��<o5�/���Z-ވ��\*��/��e�wV�xЮ)1H�0�z��LF�6)P��LN�{���@ݓ��;�_^�3+d�	�b�N��G#t9�S��o����8o����NAw�>���;���?3�LD�[�r;#��ĉ�`Y~��+�o���lF��[Hk�tss|�V������B Wl�U�*�=��^܃�>���D���$���EN����?��3�{�lg�'�G�8� 	��[�+�هKyru�	h��gF��#d�6��NɀaC�j�wU�P�TV�9�t��7��_���6$*�����P/�5������1:�<9��5�}�Iй��|���G ���D����Ҟ/Y���揪�mxF�'�X�q7��>(��d��-zټL�oAw�f��	An������>EVm)�=�c���u��~;��U��6�C�I��E,�Y�J
s4#���
}�D��wW�'�9z-�S��,�z�%hQ�������Ju�k�݌jTb���M���j
-M�E~��[/�jb	qB�/s&�o�P:�nta�^L��C��ڄ�醗�b���N�&E�
�1�~�v�^���7��I��A����dP�;����Hy��a�f�C�i?ƫs�8��K�xM�mm��R���dzE�T/� ���-̷�(C��!6~`\�[�Qa~M���.;更�@����/�y�/���{[Y�i�5��,��q2����{Cw�VTif�5������"Mi�W#��.9�ɞ�+TƝD��H^������T�m����}A,��ά���x:s������0O�����˟��ߧ����gm��8� �S�~!f�L��X���S1ax�Ϳ�P ��{^���q��cilHA�帖?#�!ݴ���,秺ѝ�}"pwN�Gǖ ;?-:gj�<e:� g:RRA��_��4�"��0�|AC)�M�Z.bK����5X@�v>1/F������{�N�l�r/�p@�.rc>��K,)�ł��g�(��幦���o�ꗨF��E���㑢�O$&L�e��6d�\Xu�F�V�~��\��I��������|�����.{���F���n����W��6�2�8���Xg[��/4@sHIT	��������0�#?���FVc*)�?ɚ
k��J�Ú�D�,���$9��/���0#t �+�
s�����ִ�Y0b׃,�Cg��`�s����,Z�d���+��v�8뺰�9nf�A�ڌM�>갋Y���r��X�޿��5���ig��i���\BB���oԉI����ne �k�z�;g���p4�i�t�f���U�F&*A�{*40���)`�'f=,/�Z����i�6�R>�+۝�J����·�2׮�H�����BC��ht<l
�m)���D��2r��WggS��м���|���щ^n��[?�D���8�a��M�@�C�y�Uǽ�3 ��61�¨��e	s�|}8S��BMz`��|���JG�x�y�Mމ뉓J��Ĵ�����*^��^|�8'bj�Kǫ��D�@`�6�h��*Z�sհC�Tid�9i�=�	�Ki\7�/2**�nX���X�nu2y����>��w�Zm�2Q�f��T�ה�D�8A�W��E���rK+�<R�jHf�{2q�ˆ���ɽEGܨ��hQ��h^k��%hۇӳ<K.�^R���b����L���[7o(��X�Q���XJۍ{p��������~6d_q��v+PxdѹLO�)G^�ń�-,��f52z��p��3ƀG�)�X(�.E�iI�%��Or�n��@ȢR�3�(���$���{�Bu�M�$i�A�+k�R*�1�����V��1�� ���.�[<�gɸ�!�8p"�ӧ(؋^#i� t�a��ʞN�8�z���	8O!K�f_ NF�S7-:�G������B����ƿ�\���]�!���U�&�kXռrsQg�W���5<4|���Ɨ��8��,N�?�K��_�7P��P�,6�=�n�T��ZDD�(��kɜ�sQTCS�EW�����p� me�&>=R���Ta�!G�/	�l�ߜ����1ʰ�r� hRF�˥q@6��d�ځ�k!TQC�mў�fc|pZ�=u&MF8�4��˟&���Bc�����L���z�Šl;/�2N/�6*�F����G܈����~����D���Wn|�s0�|�Ҙ�(��O��7�@ZSf����Uk��ĽtTWq��.ͺ��`^C*vX�����e��s��=�^]?�8�peSs����v�7�����"�C@����F~c9��ُ2��c��Ws����������9�_2f���z 
�XK`˄��4�sE iY] ��o�Aܾ!���5�i���<���V���Vd}�Q(�:����o_�t	�������*�ߓ����8��!�a��w �oZ�$�d��ׯ65q��;�n��Y{���2����W$�_N����>1| ������?�ai�F���Jc^2H��)�X$a�5f�hޡ�я�G(�Ү[x�6�`�΍����	��c���H���N{(�f�S�����wz��'�WzO�]t_Xt��*`>�ǈ*C�T-௟�
���]R�ɐD?� �n]�p�"�C-�v|{-.�ǁ%R�\e4�~�I[%��5� M&���-ͬj�i���6+����=�3�̨�
~�p��+V|v��ٌ_��`�7�Բa��B�wK*������������{N#/�fQZ��y���]l��i������?F(KQ9oFDͰ4c�h�
����,$��<7�!�	s�F�����LK\t�r�X����bم$4cF�x>���k7�Lc�d��u��{#�*�$�/6V��T����[���?qub�,�2��a!G��w��Q��\!Ի��rE��{�L��騐�/ u!���I��E�O������m�Z�x��R[�n�M���Ɋg�GZ�t��Q�F��C��-q�C/f�'݄�5��PW�Tz�.�,ݤ^)�����@Ӛ�t����}gu��WWa���_�}@b��+�����w�1w��]��Nl'��{�%���3��?��n3�@��Z�3m'L�J�L[�@!+�9�wN?殙弯/���%��� 5$�� �֤:��&�lacRԔW庉��$�&'(�D�$���4/�+�bp��s:ɷ�@�i������HP� B���:���-�'RgWd��	��a����hS�-����W��.'>�l����nإ�B�1�v;%g�`@�c4�d�4�|3����J���N�3#<�*�u�����"�/H)p���)���#D)	���c�� B�z��N�����76��nA�

G���V>9�ri�'&��w��b��^�������ٍ�űw���#&ū'� ��ֺ�,m�R�O��/�,* �v'��5,��q��L�b���`a�TT�X�5��O'z��B]�?����pɀ^��So��O�������{Z��oQ�`��˭�)�r��_oD������i5����K��)�d�~鬺S�n.뮋oz�����uV��m�ܻ�H.����E�h�v�Ն�) �Z ��))�5�҂K��O'çdd-��Sى�>�����ҵ�X�?2���2�x��dCf���T�m�0�tr+du��e�Kx�sE�1y�~��_i!��ܢ^���nV��AVe5�\���αT������>�7]hz����F*&���;6	{|�����~z�úut��o�$�$�Q^=�a�d�f���C�5���im��5��mf�/@��T�y��ڼ�1�Mi�1i�j�8m��qB�;w�푀��y����T�6� �
DwQ�G"~X=�r�� ����X����7[����;��y	`,�����>�K��*����a�A$�bZr�Ӑ�Ҋ�ڡ"�����������^�)/��U�O�Sv<7���+�i��J�����̥�*%�|K��B(w%^��Xڡլ�.I� �귞��?�Ϣ��#��i´}��ٍ�c�H��VA]<��<f�͵�vvݗ��A+	����`J�,xl�n� 
ڧ>���6�ή>�^"��Rm�难�D�]�DO&����?w�v��:`��'9��JT�qǷ���@]��P�= �%��l���ʨ6��J>�S������RoXk��:��q�o�&�5�������$v���ysQE�ճ�E:eV쇇��v/�L������aRK;@$0$W����#���\5r�w�-8)��d�#�ʰ+C���&������cB7�|�b ��ͶV�����2~�i���H˨��ӻgyƵ��K͓/Bw�A4��p�C��Fm$Q�x�4�C��
� ?48ި@ܲ�N��Cm-�/4��H�Z�⃌d�A&Oc��]���ϙR�՘�4� �?ѭ�l߇l�*�n�_��=`��^2�<�F%��^��pHl N`���?��x�W�|�"�z
��"��{̄�W�р�+��PU*�P�a�N���GM�ĥD�H�S��JL�%rܯ��3�6�3�]�"���f���[���Ia|@��5���9�(�W]���W��a�]�%ގ��a/�D2wR@�Y�-Yo��q5�} �UO�?�.�>�	3�
�/q�����u�7Av��*/�Nߟuq�DYz�(n +.�~1�"�$��%���t�,DL��W
�CaL]׼�����w'����n�]C���8�N(N���\���t3fg@�[WJ�U�A��G�
��s�����E��'0ݬ��9�(	�I�>��6}���$#�ۅ�볝#�E5Od�n|P�#Ā�U�5B��U����40t"����FDE�B���`�A|���.C!���.�j��j���$�D�z=np���I��W##�<��NɃ�������{�
�ÿ�*��Lv����&���s�4U�T�L�NN����@���_L�YX�l�!�j�]�@� �������1�h�L�ZӄG�fb��3�b�=_	�6����>d!��4|�Bʆ��")�uWC�o�C��"z˶�F^=�S*����9���]�,�	�lU5�-)�I���ewaӞ���v\_��{�HbJ�[7�٪��/�_(����\��tnW�,��'I����r�2�R��FIb�[a�2]3=���f��&�T���U�151�OgvR�-A>�X�aׅ|}2��σf�Dq�(1X�t���ye������J�rܹ��O3�j�p���R?';yՑ�I�1{F�	�=��<�F;�S�
N��|W|�{��
ʷU���Q$*cyВ��m��S��w±1��}� L�<D�@��lz�7��+u��)��� �f�.�hnt�b�\���*˹���YwN���f#�#�� �sI���r������)/��(�_R/q�<�k�x���u)�p��V{�:JZC�w����'�߃��5�8)i`/uRr�#u~S����HL�g�Ym!ĀiDh��>/���
��ݮ
��fԾu站߅���ـ۸�]n��-5��y����>���m�b�x��>b^�y���Q�A���%�y֗�?u�̰u�l.�����v��B�WC��o�ԗ��c��,��zCE_~협������zuDV��ۢ�Ę���ۉT-����~�k����Ëm�[�E], J����Zy��w4�w8��NH�V'B�����=�a��x�*��7wL��T����ؖ�c}!������|Ҳ[�7@r��/���d���S����y�1%�9&�����]�-$r������,�F4���vn�.K(�%�!��p�ń�zW���0sr[ۛA�S=7H���V�S�f�FK��6�ș\
X
��Q��Cm�ՐV��:4��A�'��o"���C(�&N.��ur����)�c1�Мp�"T�v	�J��!׍��������	�hS�'7�8�]�E:�s�ےd��U�ܨUU��[
T���9�s�I�5Uk\�f���3 �	T%��%u��7����i#�}K���)��"�Ģ���X  :[��QVݒp�[����MK����RtJ^�|�R1^Go�a�&����P�iR�8}��+=�T�'�i�]-��.��gc���*�f<��s��.��q�t!����v�3��Z�7(����~&�X���4v��$P�h��4�:^yy��m����%����0yrN^�&�d摔��|;��r�@��{@�ǔ�6����a���	�����E����;������-������i�M�
U�U��sꢮ`C:��<zi�O��c�le'�ڸ,��������aҞ?:f�{q8�%-_��C,M?%�W\v*��1T��K��@�"����%�+4i���>�h06Շ�[����F������cv�^]-#[�!/�Ř�3ۄwʄq �e�դ�G�f���A�kbk�x�u���0���B-��7'�r5��hC䗻b��-�@�>s� 7�u�_'�S*�S>�����]���a��R({u���M�Dv�"�׫�������|@)R"$��e��=��Rʹݒ���L��H�����	��"�:B��f�b��Y�Q8�Ĺ{��� 9�>
�H7����FFj"�It�<B~��Y0O���	����$�!��w�x����*�fGG�&���;J�~�5v����5��P������[�0���ѵ�b?��YZ�m���B��*�dÂ:)��<	���
ql�b����oB�u��◯v �p����x�f�/(�`�]�4Ҕ��,i�y��(~�,8E��gY.����Y��%.�|H��z��T�6C��
dB��U�2�TcjC��"�V�K[��D&�H�H��<=B6�����c{15bw��.5���t�U�:����-<a J����t���j�RB�����4%X:�w���*�b��9V2��G'��FP��φ���.t%u����+!j���
vS�-����$��%�L�@?��:���M��t���9��rEDx���<�@ P�k������% 4o��§	�^�]Z�����_򩄜1��d��|9)Xâ�;o���5�����a<=ea�G�mC�x��$?Zf32���'NF�{���ɰ6�YW�jZ~D��(
Q�����U05ƫ�/ԇ�t�����z�_�r��X^�8��q�U`����0��m᣷\p��?�T��$t���|�H�6��Habb��1p�����M��\��c�����y!K�	����H�q�+]�y��DE
�{.
�wꚙd�ũ���(5nXz["�Ccϻ�"'����.ě�`��6nZ�i����W��F*jH� ����� 3	V���c����6r�˥ݺ-"x���B1���Ol�n���.H��p!�Ͽww���-Lǝ�B�h�Ξ�>h����.��4P�r�מ;��j�s���O�&,�U��=C�.��hd܈Ω��2*�H�7� �[dbG�gl݇Ƚe����Gz˅*���`�x�;�wg�9VP*`:�|�^�Ǳ��2����9=���:����dwk�d��5
�:=!��ձ--���ҥ" aO�Å%����ٟ�����@�E����`(d[���2,-)4���ey�G�-%�i_6���H���n�7B/&ah����l�i�qk�:����iw������K�K�x?�:c�Ȉ�Ly���YeZDe��Y���I?�tA.T�27�Ǫ��,�C1�0=D�F����u-���I��)����`seٞ�H~��v��E�)��.̿�[<�!W�[1��f+E��0U��⵫?5e|U��+{�hK.��)�k����]�)��N~uݍ�f�'�����|qe )��$D�Z�7��/��N�4�#X�v�t��4 C�l��SG����
�Κ�-�0]l�դs��~��&�%�L_iƹ|�H:oy%Ҷ�L��]�E���q��dQ�5{j��$�-P�`#LIMo�@�:~�
立!���B�~_U�e�6��Z(W����m"Ђ�|��������O�����Ajq;��)5z3��W\��X3��H�7j�`'�%(�}�v3��\�A9��H�%�D��@�֬�򰑻T<y��(���T��d8��$e[��3!�z �����=M����w��p�fϭ~�^�3&=2PP�_}V�A�7~�Ӄ)SG8FO�y����y�	t���/	�S}u�8c�j'2��QH���R?m�&1}��7�C�w���S@�A E�Uns���<�p@�ҩ!z�B���k-�/����C潗��0��U�\I��\���RgH�ś^7�������b�d�����2���\u6G��?]����n`�g���: �H�	B��ָ��'�7� ��1x�ٯ�.�0]_6WD�$6���Y#�4��3Rj7Ѩ���uܜ���ҏ:B`&����	&
v��]�P��@��Ʈ�`�m��E�`�^*�D����r
a:��ת��q����y�R��F'1cyk0/K��5NϘ{0.5��V�Z��l����Я�A���-b��m�늟�&Eʽ�ל��y�RG����j�C����E�^qi#i.s[��r�Y�N$K
�}���d��&d11��z��.�0�}���K7���(SL�Õ}z���{M��y�a�����o�%C�79[8��kb��ٸ����S���cs~�
��>053ݴc�p��5���H$V����{�eׇ��2ZE<�I"	�Ư��7�Y����[�f�D��9��-��ôH�E��5^ʪ��~�/uش�l�n(^- �d&�SȬL:�t�(f/A�z����k�ڼ��?��l�'�b+�I	���H=߭�a�.f�a���[�ӿ�έTa�~�5Q�� qM:u�jB��������ޕ7���%��q�QB�E�* �!�5�WQ��[�A|��
ez�u��L��� d���V؆�&��`1@B�Y��uQ��L�C�#��p*���.D �sl}�ɲ�ţ�k��.]i>%��A�Q����S2M�*���X���ݚn��Zp�H�f��Ve�J�A��X�}�XoY���N��Mɷf��ӷ�����E�R�'m�Se�M&0��Q]�2͈��vY�9p{�!y��\0���1ҋ�,��L�p
N:k���0�mF���Q&#L�<�����,���#j��?�O�ܛ��+Yқ�A����@�}�P[�ʣ���y梭 ��ۮ��u[��6���8�Œ�2�T�7���c���}n6�����%�x�̉u`�\䡻f/pl7n��&S����y�46�Q�"VE�Է����DO�����[�1~�
(���$yC1�[�ujMi,���WQs���0��!8�}����@R���2ZC��r��X�X��5�.h�ѱ��b��},}���q���Æ>�ͥYmMr�5b�ڛ�u�MQ��1A$�4f��C��^1l��u����[.��b����TD����U�����w��;�J�>�K]��D_�v�[yCo���`�2=�$�3<�ѫ'���5�U�R��]���#m�.j��`02|��~h{����t��\Ϊm\]gft?N[\T��Nz��<�-@ͤPp���5��z��XZ�B�1Z��/�5�\;UN����s��c&`�k_G�v�;o���ɧ���w���O>b%�.�`��2长v�M��}���_~)�TlM4��C�S�K戱�ˠ<�E)�TC�%��G��mZA[.�y����.���F�à5�y�lf����Q�&� 1�2��X���N�}����^� 1��F����:v,Ej���<]9�K�{���z>*�6�ַJ5���* ��d�Pj�;6��miܨ��IRJu��3䋟sw񴤙N��*;n��O<6��<�ѧ�����6���y#�r�oӆ���I�$�Ԍ�Ї�F�_�C~��<���/�`M���vtP1��u(z���|�AWt�_<�D�&�T�=`�=?��wu�����V*4v��؏')�������P��Tꇜaw��>BZ��u��*��u��a�=�d������hH2�Q����!B&�Z¾����دok�?=}�4&i}f�[4E(�y�Wv�@#Z��:�����[���T��^˸>+0d3�{~fME�Q��JQ���h9�0����-u���Q�B�=}�Ǫ���{�m���捰g����4qd�x�t�� ��9����,^�}B{0	�]���_W
�Gp]3M֪
�l,�uh��f{w �=��ƄԀ	b=E��f5T(&�R�̯6ҽ
N�dr�Y3:̅4��&\�
��A��e׃��S�݃� Xޙ�l��ȼ�TM�{��)���W���a:^@i��g&�g�	kJE�{�i��+l�m��bk�l���)4�~�������kV��»-���_���ʵ�eJk �����4�O��17Q:�ȉ��t��b���`�8T���v�����?��K����´��N�
���8g
��+d&�<�x���NW73�}�0�_}���Vߗ?��R��4{s@)�ɬ�׺
���p\�zO���;MPQZ�6^�D㚁w��RVd�tC�u�CP�@{��O���`O�UaQ�,����	�D���W��:��� �8��E걭v�rY�)�;��A�Z��)��:�C[���S�j����Xݜ��������Wn[Rr&������'3qF'��O���V����)ĩ�t��h�- 0���Ӱ�������t�B�8hJ@�@5N�ɔ�x�p]�g/���0gƔmG�O�w$�C�h�P!E����'9o !��2w[�����5������,eI��u�C�2�,�Ex�Ty��%���9m�ߗ3��Z���`$L1!
�h(-���wK�I��/@�y޷�Qm��R�H�=��Ie� ���f�������FV��.����D¾�_�#)`�An2��]������1�@�mN8���9n�w�����q��G���|<���G�1hN ��=6ֳ�:�r3�iE��\���a���P�������(������l�C���ޕ`�Fz��)q�y�J7[�a;�g�i"�ƗO��f�z���0'H-{���������_E/���(����L�>��N-��`��������lǔ��Ųi�l��S�͡��|���T �IQUNaտ8��e�L����G7�zb��_��)��LU�S:{��X��g�vW��_�`��@�ﰒ8@�t�P��Qk@aeh՛���/��FYG^l3fN9�ۿT&�+�t�Z�h�^W.�f�;�VH�
G ���}ܱK��޳9s0��J�J�LP�`O��>	���?}]�Ĭ�L��g�$�_�A΍B�2�8Ft~@��I�j�wy���Nl�U,p9�zZ
�m/��~��.+8�X�_�D��KK0�u��,��V���;���T��mS<�y=X�rn��zuS�J��<�ם��uJ.�jh�����4��As?{�c}�`Pa]���I&.����7�e��Sv��j����a�}H����,.��4��Ѳ(ּz�w�>��⸀Sk�˝e����Dp��M)!��b���6_�lp���P.��1s����=�"\~���<�l�{��ίz��C�^�p��}��bC��roKL��Ԡ�AT���!�������V��m*N�)AV��B�ّ�����
����8�1��L��]�Bm�0I�RJ�H{6;�#��g�1�+��G��P�q���	�%y=��f��!�vg�7���w{�� x�0��;�]6rW2�|ڿɷYSG���j3�q�������L��Kx'��5�V)���7��~�EV0��g#�rRCRr����72���C��T��P��n�ͯ�Gh`6�����OU'��߯4v9W�u?TU�u4G�{�|�g�v��ylp1��R�
���'��<���T��c3R@X>n��DewP�v��QIV�_T�����Ww+>�V�谟i�h���m��oǁ ����8XXdSl��S���,��SkДN��K��V�Wc�O� �@�M��D�<t}6���8 }���nA����>���4��/�^�E6��ݝp�����<ɹ�/5��"!���vw��ҏB�������qS�~u(]
CU|��ou�)�m����@fm+W,x�NL��%iH8�T3o�K�&�޳����\f�D۷`�a>+�gH���i�z�t�$F���QY�7S��w�DÒ��&o�Y$�u���]������1��+�����[���u�U�=h��	���jhYr'��U� Z��y���ۭ�;0�#l<�K�Q���w.�MHP�v�J��p��8���u8����2�QE�z
�����D�'�N/�k�#bA�ђ3��9�uᮠ,�P���wh�q����2��⡀�� �e�,�]b�Y)X�yXy��d=�ز�)pwB�]�X�	AXl���f�M(f9��׹���.��U(L�5�Y���M�ޚ7v:��YC`���5����¤�j�E�1)\���g��"�p��{��=���+wWcR�Q�M��/��ފhp#ե�j� F�5!���N�G�����YCAh��ҽ%��%>�Z�Bޠ�2r�߻���wL;���m4
�{�A��7^��2��r8N�7jj"�O�-!�ݗ4nj�k�m��4�����0'��?��p��O4�����6��8���A�;C�����6D!�&8H�q֟SdH%�{6
Н�_]�
Z_B~��_��ó��Ch� 5MH���a��$B�O,���R�N�N	����<�8�ղ�2�v�x1��f�`vN������Ʃ޽Y91҃��q`��Jch/��w0�ѹ�1��.���/G�5�N۴+�ث�/���`�/�NS�B���ۤ�Z˙8v�^��[,�6�bIg���%�1�����9�����J0�%�ӏ�۠T��=B��4�p���GR��ð�א=ci�ˮ$��c��IH�[���UX�^x��x�7 �)E<4!M��x��(��2�H�y%��g��������Ih8�'^ Z��h�^+��=)���iÃی��q�������{� �\�M���n$�X %Ñ�7�PG�.�3���!�h�FM�fty��?K�8�g�>[��2(c�K�o�+ζI��v���SXS��Ǵ@I��A�U6#��4�Dz���_��`@�W���35컲�P�b֡�ӕ��%L��5	"�� ��6�ƫ� 9��[r�i�-Ĝ�n)�rD��c���y\��!��BI>O��FϻD ���(b�8���8�t"�d�T���4n
Y�6蘀z,7�������b�+�p�i��Q#��G���n��hі�8!2o뺧�T������*Tf 2&��z7^0��Y7(���?�ģ����0�5�L%�F���*A�G	��]&̩`"�"�>��p�h�h_)@e9+Q�毆:z�i��f,�7��"KkY�b�z�깞A����
����κ��V�gB<�[+r�,H	��NW�2�ǵh�7S�rP�Y��������2eO(�4v�yw<d)CCJĖ���"��Af	�1�U䙅xXrM�vȮ�$U~���q]D�g�G[�&k������1 -�~��yO�������G�� �n���Q-��'��#mWS��a�ӕ�$W\��B:�������*��~��R���uә��-as��6
=�5�ג��l��*jU�MR�+��;�1q!먾Q����m���y�4�<,��:cP� N<r�3�~v��Isa�͚&T��OM��IJb�G�5��X�c�O(:�^ɹ��+��:a<ʘ9����J����� ]9ѺUp� �M�.��/!�V� rT�sGt�x�����{��-�Qٵ~�n;��A����鎼L��\1`�
aOWQsX\��-ʿ��Q��Gb��q��SKxG���#_�F���ӊ͗�&���Z���0��<;�@�'�x%>��5F@G�+���m~��Z3Y�k�LZ�h�)�x���
�j����dc�}~�G���C�C���}���Ydq)������5�����I.J6b��~H]�r^��#v�cbs�8�g,]6;�)��q��������AM���}��[�M��WyȬ+@��X4�;0 5(�>l��(x�8I� ��f{���
�-�����"��Iam<��`�Uw�0"��	n1����Yk�e����|߅��}�����'������3�!����=[ɫ��#�����[�)�&ԊV�� ��4O=��ؠj�W�'��8[��le��׸u��ߒ��[[ж�D@~�6�PbU����F�G�J6��> ����)Z8.��!	�N�A�s&�WQ�|�Z7s<(ܮK���ƭ��d�〿UA�ݻ�s��K�pk��SFP�2��bUK\R��[���F����8N9ª��5��X ��(T��$��'!�����O���6zN�P9։���K��CƄm_\�z����].�m���)�j�C�f���Äͼ��b���<_d�Ժ�H�XN��8������9��H:��EJ|��d
��s�g|8X��	�U���Nz�J%�����`ϒ�<�d�G��̒f(Y&!�|�&���-��6[\��9�0���o��FupK��G�o3���^Q�mF�o�qъ'���I�)�4 �0�{d�_�\�dPޫ�tw��:�=}<�c���!Lt=�~�.���Svo�I���t���_ݯA5_U���`��7-��1#�n8yďa4!zE�B�HMxW��9�j��	�-��BN���d|�3�WQ.��s�O|�g�a���o����ʛ�M�ط]�Ka>�H9-����H;�9~�h���
L6j�t�:���v?��EI0`���/ͪP�\ͳ�8Z���Qc�ެ���������W`E���0!u�7�ޣa�E�I��EsY+���G���nX$��l�)\z+I<���\%��F[��~�q�45Z�Y��8�iԆ�A����"�!
7Ir�=��rKv�v��g?�G}7����XH����5��Āw����.%��{�0̘���q�fN��G�F<:+�:�R&y$�r�����*Ã�)+�/����yqބH�d#�q����X_H��Yi��Ʋ���.摇k�*�e�v��Q�rG�t�ٙ���;�>���fI�j�����F���&������Q�g��J��J��ҋ}.�G���2�I<�aس�8�}A/�K��1�^����K�OY����I?���oIK���~�u%�T����iDr^�6CmH�G�#s���mf�Z�,�, ��:� ��q��I�b�`�����|��i8�;�!�R�}@���갆�r�G�NV��`�)+�m��(S��ª��`~��.V�=��A�GVʪ7&򐪓;��3X8l�ۮ�F����c�c�f4�	;8�k�.�y�,l�P���Y��{���,�!�`���ii@y0�6�)$}3��`�Z�><d�q�Z�c�*�e�p{���WW��u�.�f=����!H0ۭ�p��{�~I(������t�(��{�$j`|sa��L�})+��2x2"w[��U|y�O��QǼf{<l��)�z�U"V8s2I����X���ӣ��Po�Nי7E�M�������՚W��hU�t�ӺV��?��(�>����oa@�m��Do�2<1KN{��-���^bk�x�����v\��Ӭh����a�v!�{�X��(�itЭ��aEtR"�	+'Ȩ�sw¿RO/KS"!H0��C��a���&o�C�� %gM����!Cbh5i�e�Ԓ��0
���΄��Dq��kk��D6teȫK1��E��C(H�*���@ʛa���*��<�����|�a� �,���.�{�d�pS0S���lN�~fQ�g�9N?DB����� ~LA�֣U�/�-�8Oc�Q��7t��r���lQ����M��X��K�������<���Aѽ��l��Bo�6\E��J����W���[���?��:ZV��Y�'���.D��~���~���$q�����lUa��C/���p3�p�~80�����[�#�i��w�%�����E��Y��Nc��ǻ�3�;Gm��7Dr����Z��I��]�@�x��������!��Jcw�NI��F��-l��&=��d�<���&�..m���,���.������7��!f�˦}��;iMt����2�yo��Zr��7H�\�6�;Q�����+D7h�(�{��(vh�$)ش��Tծ7X��>D%����<�i�ƚ�irwN�.E|�5fE�@7�a�'��#:رL\L���c�W�L���p�P��T9�Mo�i����_˹�*��Rk-���:��N�*+�_R�^�[0m���#� �7�w���*{�|�)ϧ�-�Vj�z�]d���+��8����d�p��︁Ay�+p�[_8�����` F:�s��m�a���>��s�!�|����yª;�W�ElAb=�⟚�=6��h	�����@��}F)_&���e�>�ψ��EEy�W9.���m�%�䥀}2?A}l�{L&��0klc���F���on�B���}�+T��8�1�y���&�
�K����~�i{��tl`Q	nr��B�2��$Nm8�	H\?.�Ga[��4�lj0�O9V]7Z'T'v��Ic��_�3)��l������%��4<O|O;�~��Ͽ'c��O�#��?2P ���$ו���%��e�K��7(h������d�s�"� =0m5�,b�;�]��DG|F����D��$�j?<�*1�Ì��g~�!�%<�]�	�u�2O�:���O�BU�~/�e3.]��^���P*h��h��M_�er����x��9
~�jQ��W�mml�yo��i��ɸ��	�椴QP��~-���/ú�SsZV�R@�'ى\�x(� Qt��Kh3l���Lr�V�[5�#[���RHK ]0M����ln'�(-}���JZ8�-��*�-:�	�+�+l�����sj���)�?����*Y�����)�Ԍpf��G
yq݉�I�E��KP� �9V������ݩ �%�6���/�d%���XW�����o�V��'0^��H��*�,cٻ5�H�̙{��c@���9�]Kos읒%�H�!��mb),Q�s�\_YǡS����6g*z���> �t6sT� f���ʌp�f�2=��7��M��B�ۍw"63���Y�˺4*3����UPg{�* |�\"8��쟄�ӓ�׿��N8�;��h�\cc�௙�Sv;+��tL�h�f��`�dIC���"|��8�[�'G f!��Ś1��Q��l�	��T��.^��OF��7˟{��ژ���Rxj�39��]���_�%2�HN;VLˆ+fi�D���a�T��S���#]5'���p-�Z�7�iI2`HX� �DÔ둝���*�q/�vu�{�Fʵ��p���
|�۱�0�r�,��9٣���9d�)���ld�]�<,�f�،�-��3L�9��=�&p�N���	h�d�j�J�ﴚ�;0�	<7�A��I��d�I���@�=����eH�s��x3�쫷�>��W�N(�.ᆬD�(;�~[߃�����,�<�P;�RIA��_;���ܸ�y6��g���¢}I�;��~��A�?G�O�$��ͤ�Rx�*��e3͋ :p����\�&1��`AQ�!�:S�UnC7u�i��h�ә�	�i���/������[\�Ԡ �#�<�W�Ւ�Z�y6{��U
\�V��@��/�X�cց1�sE�vxp�a!絯��E�ʐ��F �k<�?W�^� %��q�M��- ΃4���9a!�w��.D�ɰE�V��ɢ�Fq�,��u-��,��k!��MbM�P��}�K�
��#7V������d�JR\/�~�)+T�#p���a�#��0�#m����v���2W�������zg��1��Ч��Ė�a�����r�F�ֳ�L[���BD��Ǣ�'���F{���TGŌs�w܀aЍh3�ͩ����*O�X[�il����BfAV��`�g?Q��.�{��ϑr-(��s�����o�Y�c�$��oU46��C. �_�X/��ZOۮ(����q �h�����~lTh
�����˼tZ�/�t���!��?����%�[ȁX��2�.�����#^���t�4�پ���_�Ͳ�\x�u"��q��xJ�L_L�Y��f 9L������l �����񇎻Q4�|���Ց�=�{ fJ��_R�[{7eR��I�܊M
��Ow��J'���iӼU��v�Qm�����%ta$F���j�r<8PӖ�+�ţ�����R�]�ӑhC��J�@���m5�����ֆ���5��C��G��,[�00x���+�B&��y���������x�B�x2��NF>�T��YI��ls��ĕ�s���R@V��K5#��(��g����e�eؙ�_G�p� ���*��E$^�8C��ڐj��L?�xg����r̢����i�~��!�U���wx+�F���¥��|�S?���_�'��o֛3*�}Vj�������E�ٌ_:J�c4������J�f���X}�AR^�F۶��Ľ	��'zN��}\�����[Z�i��h��d�3 ��Կhi��H ��x WB�ޞ�ij5��K �h�]���WN����"=�F����fA��eh�7�o��w�������	��w�W~t�#	wl�6��a������/�H��v�
E��W�Ԁ�*�t7Z�&�B~-�EH�����|z���UU��4���J���M�E%��h��Y��~�tL�{�6{��kϞx͌�$Y��  �e��p����C'b���uZ�ND�丫X�J� 'xW������_�i��U�
�yU]Dj�c#:�D2vX�:p��<�'�}�vh��,/���ʱ�ZK��ŀo6��
4�$A�'B-Im���E�M��Ի���ߍ��%\r�V���"�
����&Z.H���T~T$��;����}�����B�M�����������r�y���«\��q�=t��̈F�<����0L���Dt��>�1~c��t�v6?9'� L���B��d�~o�&Rhh��{�=���8�=�hd���BD���NR�c�,���[G�c ���O�Uz ��O�oe���p��M�N�U|�^��@� 1�͇��8<�����ƶ�����z��'Gb0e�ά��9SU91��N�B\c|��h�Q��W����AT�� �n�n��[D��̵<�0
2�"�D|D+�G�Gõk+�w1��F��+��Ѳym��=���j��<J�������K��0�\��ݲG��t"��1��[��tX򗾭L�)k��|����ʌ=q��rxM��c:Ԯľ�[����m��1�1��aɈ�&�̉�0���z�*7��K˧{�T��Y�؎�$�����K�]�ø=�_\~�}��=7�s(���h��C��e�bq�FN��%�+v�㟑TYFU�J��5>!6Ř��T!V����&�#4d���!@���G�ڈ^�����垜��0@&��4�Ê<� xi��_)�;��A"��ˍ�~�sid�.��T��DŅ3K��a3��♔f����1vZ#B)2�c�=:2��`\`Wt��+�:?>�;Ov���P�d�̤���i3�4���!A�4R����`?Q����6f��5�oñ��e��ꘄ�������?��*5��x��,����j���`�(�º�;-�
�<�4g�JR�rw�G@��jm&�*�!\	L�ʩ�rz�� TB�F8��`��f�(�UTg������hE��q�m�[MWc��6 U�	"��ϝ��5��`7���?�����g4�����)��d ���P��#�0�c��*��y���Z�n���c�pRH3�ӕ��aUTq-�����7��n��~C\����3"`7�B�ub�`�[����l�DI�k؄�;�k���9���G~e;���\���i�:}��}ʭ��)�7����2��0��	�W�e��I�Go��H>����J�m6�b�aJ0�^��g�~隋ۛO����ɇ�q��@�:�v�����ICѽ7���E�{��4��\�
:���b2��2z6c�|�WH��F�Շq&/����@�d~UI,07���� �L�q��ˀ�J_��pNI)���]����}h$��⯱%궀���r����00Pp,�8�b��z3��i�yGˣ��Bo6��)Pi�I�c�ǿ�"�pT��-\n(m\��w⺟������\��%�e�V��(�y�9]�Ο�T/�R�D&�����X�����F�S��D��c�o�(ޝ����=�JY���/j��%�#NO �2�, �~@S�P�m���x9�٥~-J-����z'ҢPq�Gۅ�$�\�ICIFN��DB����]q+�K��t
 J�7ւ��k`�@D�A3��7Ҩ*���}�{��!kT�I�&��F#��_9\m	��s�@A�k-�*e�C|�Ɠ�9�|D��h�а>�v�s*p=����B�T��W*Q�%�����ߣ+���3����#0�x&Z�Yű]�_a�ϲö�ҭxȜ+�Ҵ�v�<�����1���T���!����%t��ط�����'5��4dŜٱ��D�P7���qQ��	��!�SCY9!<���PE��]�E�ILO�K���
��@�� ���ir�iTܥt��H�R�?č��Ө��v*�� �\�7�D�6��w��Ie.F.�	p��U��=7p�����v:��mwu#�0��O�O_쇴�s���sҷ��1�yi[��D%F�2Z�@�H:�"��qOW�7�J�.d���:I�dMtщII�j��P�teЦ}�����	�O\�bK,��DC���_�d�n�լ���m�0�tZ*�7�n�E9�6��'К�hUt����o<ݒ��Gj�~v��{�ͦJ!#R$HA�M�@tc��������%zxA��V�Ԯ������U���w��B�N�Zg@��S%�o��lz�⍿��;0J��R����$�z\�έ����w%���>�J3�U�Bt��?��m���R4�WՅ �]�p���;l���zZ���H3�1�?B��{��t*_�n�,vF�Z����q�|�Ln��.�(���r�>��"�v�� {sc��`,�P��挣 �4�[3b(W��q�m�]���-���TKSR������+����V>SNs��u�ݭ�mr��a)�,���`��^�vhEsCb�E1S��ن��%����o0K��.�V(��X)3l�؂����#�|�?�	4v�$���� �������-7z���>Q����Lg�#�.s�d�Y�Կ��h� ���}��U8�\	D(�,�U��S1~���<�41�;ѹ$-��I����ƙ���o����w݆C��,��A��� �0T��d=n��R�tz�ی0Z�3��9��X+�-Ӳn�������LT�l�0@ﴚ؝�P-r�%��[D�K�?��>�nOr��5�!���-GYg35樕�@>���o�����cT�R�x$1@�$��$|}�XI+]X�t7f�6�	d�� �e���A��}�*�2�5Gr�]\�@Pk7;��l"�W\c��ф�J9DyU ��G���1-��*�%/lDT��EM�W˱��_�qY\�ty���!2E�����_K�*����Pdyv;ʙ	�'W��š[�j�c��2�G0��'�8d�I82:-�yf��n����ŠRdￋ�����d�������I�3���W�S��2Ϳ�F�%�/�BUJ��yދ.g5fcƜm$�^���z�yk7%�'�@<��9T:�-#��Z�2ۀ;����6Yh�d�ZB'mU��0�zik��#��$@�Xƥ �c$=���iį��%�£��/�l���	ƃ��v����i�ږ��s���T@hV������b� 7�չL��@��`I&��s�`���z)����`��X�m�[-lˤ�R�t?�����g2T��Ə��GSx���5g���M]#q��TvO��7���le��(�)����/1���-�C�1h�hg�'�9�(�,uj��,(�&��
��H��xS��TK���I���=@�e-]N���W
���tTيȎ��7�f'�(���Ҟ����<��^wT'>�E��L�(j�������#����RE�x����0��ΌZ���^�3�i� �i���>B��X��z^�T���UQV��v�����Uv���WR�{� �<����g[��l�@��J� X��.2���2��ax�)D\�����䑬[�Z.!�5�@�H�����a61EhC�.��ZuB��F���.U�o)�`�[]�଒U�ŃB��ւ���y8��!@M��9 ��V�(��[�C�=�+핓فy�!��ֱ�R���y��DhZ�r�T�=>$�7�5%���6��R�4&'�� s�k���<1c�;��	��g��Q�jf��F����$��m�������"Q���hB.yv3m
��Eӄ�	��x�;�a��G�5ԍPb��[�96I;C��̿`'$=0HO��[:���VI/�oB4�cЏ�&�.)Ҁmk;Pi�W_�Q��9ɶ����{����-&h17}v�r>��At����{~�AZv�W�,[��e[.�AL^��~yEh����W�V���r��d�Ҳ�>l�H7�JhO[�Ӑ��ᵋO=7W�޻�q��+���q�x�hP�(!8\f�Ӻ�Tܱ���&H�G�G�}ꐼ�.�:�E�?f�r�:|��	9B-E7:r��=�~;b�����H�Wݷ�[Q?1��ľ�P\�j
l=��>d���c�5�xQ���u�ā6u����	9�]�U��>Pz+TA��ȯP���e�3%�f3�i�&q����[���q�� ��	�d+۾��	�d��V��a�fe�kfm �J/�)ye�sT�t�:�ʫJ���r�$y�1�æ�s��9�1�wE�U�� �:�Lq��F�	f����mX9�Q��k�G�8:�n�b�:�*����j���xzIv�A��|�J4���J �:�q�LX���a���L�ıB;kb�J#�t�/�>/`�H] ���\RD�<�����7ҹ�/��X�/��^J1ph$m������?d��pGk�ǎ������ �	�����i��>�`�����/���l��W��ݒ���������躬���Txb�#!�)/? �� ��B7��5�����`�D�,u�h�!�G���h����P�fC��z	���~�����ʿ�3���~ 7J�aW	�6qv^�x�cb@W~a*r�����kN�2�4��pe���dz*i��}�}�$��4��s�`�x0FRL�ZXc�vK�$��������׋̼ja��g��-���E�s�O�&)��i�K��o�~��uTe�]	W!zJ&;�81�1x��W�L��j.�)-T��t�߆�^�w̻�B��O2l���6���]��:yn7p��N�`���ͦ�w��q�a|ԡ�Z11��V�?ҷ��J)�ɝ��8!������n���+�wc;��8��U�����c��0ֳ�\ ���,��39/�@q��/���G��w׊)I�G����3O<6�֩'���PZ�4��7K�*P=�?��t��_N�K�-	\#��z��C֘��X�twr�4���:I[>�kv�拾R�}����1x=�C&:b�+�V��P,��c��X�+��{j��2	㋥��!�8Aŝ�ӵŃ��Wvc�e�?��y�<(��`Pv��A֛�cg0`O�Ϩ���n�{����{���T�A3H6a�髮 �ҫ��)EN�!�!�:�&���};���E"�V2���d��YT��l�I���BIȗ����Q��UO��I�.sb���6����g<��#����e#jP��P��I����䳙#���7�)G��3!TP��3�R��%���o��Xɂqh5�!�NB�s�@����n�EScc�Mv�K�4��������_��5�V���H�W|{ę:�	���Z�vd����=�zP�,j��H<��^Ҧxr��!�`sO��ĝn�;)�.�b�}	�1�9��ro�L����/�6&�gg���igD���h���L�ʥ!׍�"�#�F�~��������Ù$Y�k?�����L��E(�N7�!SI�9ʳ��఼W:?�k8�sq�'o�T�����j��'c��<d����:��4��
l?^�������X"�uh�1'1�9����嚏8U������<:��e��s/ڝ��EtO��(i�Z��k�m��2�ۤB���{�>��]�RI�\���,[qa�G����<��M��M�����1�L�����|��wߩZ \?2t�Mֶb��q�q:�D���^�	_ѽ�6Q��S9���2(>3��\ZH�6�;��h��2�[���aMoT��h,:�15�P�nu�&c)�X��~�ҕm C��9�f&���!�弸����4����~;�]r�a��.ZE�ȖP���"7�P�Y�#�nad�=u.�[,�:d�ÁJ��6B!�Vg��V�ϖ��ఝ,a�զ\�_�j��}Z�?m�U⛃��M��rk,~�@c��/�&0Ge-�y�(��<�<F،����J)��E 0*�S��}����ëoT��� �,�W��R�A,3]�.c���Ѯ��ソ�Q�|�s�.U1N��_��"�u��� �8q.RD`V5�򁌇�o��jO��f���З@���'+Aj�#<���*����u�fE|`�����~��n(�7:�7�J���w���'��ak�i�g�ή��1�_p^��ց[��e	 *����?O��5��Hc?'QS)���=h/:LH��q�'������1���������������]h�ѝ�[�Y+�V����.�3H;�D��1�z��*�eJ�ʪ�"db����4���zL��2q��#�=�[�W��_r4x��':�=9CS(v@MM�縇�XCQaJ��R.<[�%Ȕ�.u�P��}l���KH��c�7��-��Sb��sZ��5�,5��&��Iи��f�����n�0�� }ź8q����?ie�ϤO��g�w�R~�ߜ���� �74]��˻2�E[�c��o��U��<�zB�6ݓF��P`y��&`a�����'���s���ŉ7s�a�[�(O�.1k��D�����S�ɑЮ��SNʅ� �CUu,�ڒ[��sM��z�9s��.��/_�H2 ���\T��;�n���/�~Q?�ز�Uv�>箊��h	I��S`�IL��q7|�J먗���ohR�5���z��>�m��� �Cc3��?�t�-0d�&ܒ=�A��aOD'�b���i�ϛ��3C�2Fv��z��dx��Z�"��#f�x�^�y���Ө�f��oz����!���v��*��q��Ra,�+�L��p�{�蠯5��u�w��?�#���_r��E�kD�H�	��N'�I\�Q���|�H <��k��H;sf��ϗ��P�#~r�Y*}.�{���B�ҩ/�ww,�l*>���S��1���V,��	Gԗ�J���k�\�[[m�KSH<�/Hyp�dȡ̙d��?��b:��D����x=zdCS�&yZ�f���S�TϚ��l�L�#*����o ;��N�K����o���:of��rxb-�i�2��'MO&�ީ���Y0f�&���i���a���8rg����kH? 4��<�lW@p7�g:�#��~rl>mo�Ɇ2^���D`�����v��-UF̾���Z{�`����n.�4<����u� ��P+!9:�x�e�h�k���1)����gS%a�L���B��B�~ #����b�������`qv� ��=��P�0y�n�|{�y�L���|xg��z�͊TQO�	&��pgq��*��E��{`�-9z�]^ p�W��裇@����ɢ?�ؓ�$#���┿iݴ?4��GWC͔��~��?����%�<)���O���6F���5�0��~�=NI� 4����V/�oYh>{���ˇ��B�ǻ��tө���
�}.\7GK����Æ�O�ڧ��Nl0�H�{{˂��vP[,��6X<h�X��#�N��7��4�D�w#��*6��=2=�;ˆ
�� �P�n��Eiw�ǵ��L��$�2�ώe���%%%ﲘu����j��
���6Q�̀(-�|�H������ۣ71Eb]|����3�?Ļ\�^"Ck�@
xVL�m��#���7��>�TX��C3���Q8`Z�{\5u�+�&*f<��B�D.4­����v�wI���������u0��B3
�iE�e���￤�]a��#��vh����Piv%6&ӗݹ�K۴PJ���gk\orOK,R����!"���b�?u�פ���~��ؚ~��3�q�]c/�%�����A!�H��|�����.~�e��u���	kXۉ�߸jg=����m)���jcC�"o� yԽ�$�4�o��9bjg�ظ�|'�g�?T���7�����*����YQ1�)W�����������dz��Yx��mzS	�lĜUb̭j#��n�F�g*V`�CBw�=~Y��"�'�7]�j�m�C�h>���̭:L��h�h����^�����K��?	�~x�}�M��
�_oQ@�jeM"�0諸M�b����sXS����gI
��� �ב���銤������:�z���FDF���r(yje���_�3��tS��ӌGK���f��@���.r= �w����>��@��-D�Q-Ts�F�7@�?� �&�UM��I�� ��j��U�!0���}(eR�ʜ05kJu�@�Sg�5�K�`"�S���3�V��Y��ȿ�{�{�k
�H�������O�%��P�+�3I&�[IJs�Y!�
������N�b/Y_7�� ո�����W���:[�%��v��6AH�G��u1��U+:�K��S�%@
v��𳝄h�R8ܾ40�0��0��;��������`��n�yL[7ܶ�;lr�&{)�Z�dƵ�3�<�/kP�'C# ؕ.���:c�ef���Q���.oQ��;�ĨbLT ���cFF����N����p@��+�ex���������1��Z����mRjR���筮;����ȗ����S������/B���n����s���ت;Y�l�ɛ�w�&|���E����mtܞ@��p��[���3ra�B۵�Hdߥ�����.���H��y��#��+��{�{^%m�vd����M�sp�K��nܜw�֒Rd��/u��5+�c-+?�/(n's��}�GB�@�	���
ku��nKl^\�c�?%C[�A�e�|O'#'ºn�mz���.��RE��c�&�Ԩ�	�.-8�6��_�Ǣ�J�
�R�g\xt���Rz���}��jo�*��Y��yvG�p23�n�
�fA�)�#S���t���k��'��#v�Sb�R·e��
��I�o���s����!wM*Ƥ/~)}kl^C/�X2�W�����b,)iv��<� *����02a~h�n�%c�/��E�Y��|���3�w�������mH�ab^_�0�.���fZu��H]EeP����f��ڍȍ�\�k��G��N������XJm��Ɉ���,YIB��E
�M0��x� I=f�=��My�",zJ|.���(�����w��h/������a�5h����m������Z�P���IT�����J�c�W� ��l�'S�:Y���Yh���X��P:���B����0�N�xp#��(�M
L�_auX�K]�p�8�]�L�T˘͖�����	��7�ϵ`�<	xėf��w��nb������.�}�M��P�y"��/���l���m��v�(�h6�}p�G^euMwD����� ww��R�K��
z�*
���+����J�E��Nڥ��*� wB3h�V����eX�Q\L{cj�Q�嗊�~��gJ��qH��(UG	R�"�Ə��h�д�Z�B��>r5rԶ9�:Fy*� Zb�Fy�����S��#8U�÷ζ�!��t�7Ubф�C-w��н������r�Ktvg���;�vGϬ�-����I�&w�UD�M�f���1���.�д�S��6a��2|�zĖ�3��bO��;��x����{�8�����XR#�h�v�Ŧ�|�J���_��%�//���������m�(]�� l���ҏ�^+��S�����6-�!�@��w�3�޶�2�y����Z��$]�k�.�N�wz�V�u����7�X[^
0g!bO�&[=�l�B#4% �/�7��A��a�g������܆3ۡԧĩ�Eܕ�t�>[�V>o�A(�hp^��Ļ�����&��x�M���MS9 /�U3����p���uJEG
Y+fU{ ��<�^�����4R<�8y+2��vQ���̪ V�+�U	C\�ǎ�oM��ñ�>�*��':��c+j�h_B���R���J�۶oM�3����`�	���eX�g۲�,�����U�2y�*T
��
"�_)��@VRv�Ց��ͶEi6��Y`i`��1s�suki
}s|f�܍2j�g�I��&��ٕ��OM�� �ٜHg��z�f��G\�5��a��.R�uf�}�g�	�!�5�����ל�4"azy:Ke��n����a�����7B˥}�߅%����u�'�`���59��(?��c6')�!L�t�m�	)��a�j>�i�$2j�5M�/y�p��f����O��i�Sk�=9�GkN�1~�]J^j�'�!�Kzn���*5�N��!�6�=��(I:h���%"�iD�5�`5���k����>��D(�,?Ӌv��40@Med�.���I����$�V<,O���	��7k���q���@�J��D8-S�|�
 #��#?��	�hB��/(��W4�)��"�jJŏ���A2�ԕ�Q3��E�~��)��ܚ�0f�w`]x,1�$����Q�q2=𬜙Z^0�������#����`<YLYܞ�I^��J�h�d�b�y"�2�ذAΒ��B@����ˬ�!_�l^�b9���Q�bn�p���6F,m!N\=鼱�կ7[%>E_��j"E]B*��jc��+k�YNPE�9bN����X��C��A�n�|'n\� �<�������c���2)��t��Zc���@�,Ł3_�(0���%�WY�v�H,��EZǕ�'���K����p�����I�t���6���PE�Wǎ��!�ލ�x�._t;����9JS�dR�����h��5���UhɮX���^��w��Nt�㭣B �ۛw��,�j�"��ŭ��ۡ-�T�n~��T�L�=�
�Ii��
�F�&���-�H�Lnȿ�j:��Fh��6��؅fs���borx�z��� ����:����z��,�Ơ���"��*�vfS^�Qy`9V���hџokp��� �`�a��(!����J<���}���-w6k�z2f6$_n�5��4�cf*���q����*����`�a&#��O�[M�8��ݹn@=������6 �����ʿ��4�=c�
h!PQ3���_3�e+dT����_�ۼ)oRY���*���\��[��'���q����	��?5�7��>|[��3l���zI������?^1" ��N"��\-1x�N�H�C��Mr��>b�G����u:����ӏW�%��Fg"+�7��d���q�s�i���0cy�[m�?�7�.��i�O��(�ʈR��O8{@�+8U��� 9u$ �O'�T���oɗ��8�M��Z �'Q6S.܌�u���GMj�5Ԧ�2T�v�݇��n ���p)�D$��8�x�7qq�!��=k��!v�����ѭ�s9UC�J]�n�*o��W=���	���=�4�`����h�P��J #O5}�+��.�'Wl�)�Ej[n����}Q؂~�;�I�F�\�����=po*���K�|��7�)��q����%�7�,p%_4]1nΈn!����u�Pၺ+��y��s&��rA�J�?�54XT�!�2*�iXb��NMB��>po�5+9c��K��_wM��2hE��'�8zE'�ZR���� ��J}GW�\�0퍗B�QZn��/I�. {d�Jʸ�\qC2d8�x�!U��HN޿�E�s����ׁ�ɤ$
�q�MSצ�����6��®�p��5<��W��+�p7o��"�N����E&�K�B�k`�`/�~l��1_1�8�M�c@6L���ެ��Y���.�M6j@s��#7���U�ĶɃ���0*���6Ă������ŸĂ1�^�zA8S�7P5C���u����
̅�#�kq*"tE�:�w��z^�;�#����}����Ǎ��v�E�h�`��:YO��{Fc&���8�=�K��@�G�~Jy�"~�z6��{�`4��.�bm�q��6K������>}Vw�YK�*9�*3�g�wo��VxR9UŮS�JalP�go��uv�h��Tn���e�������2�~�/�%��a �)1c� �׌aE�qQé1�z"���Κ�7�H�߸���![�Mμ	v�6�@�%V=��q9(N��1Kz0�H��z���ԕH���w�����$�]�@���6`CF����-t ���,
d�4]<�����_r+55�0���/�||>=R��}
��D�b�o�Ɲ�T�x^��
Ԍw��4�b�7�Y짬9��#���3܆���IBJ�4�y W�쮫R��r��S4TH�a�P��%n��|����F&Q����} �Q����/%��ݓ��to =��Ix�_�Λ��э DX��`�F�9 �|@s
�zF���9H�{Ԥ�QNi)Zq�0��=Ǡ\��?+�3l��R7�+��*�`����T�bB������<tѶ����c��(g�͂am���<9G�]�����j��ԯ���/�w���k���z��N��b>M!��PX���f�8c�:<q�v9��`�|��B&jB;��kf(��I��*-4��f 1��ɪQ��\PD���.䑀Ͷ��?2�x�Nn�A��������iY���v��e9Z�B��dI�*昿8��xk��o����Pe���&>R��R&��}����̭�u������­�[�H|���	��Dh��e��k3�ؕ�-���5�TMlZ^��<C颰�N��ea��s�@�e�%�?{
�[���f��޵:sL�HQh� ��ܳ�2���U#�~�)���Į�ї����A��ߏ�?\�N�C��{���R�6������,&�1�*���P��|5n.CU�F�K	�'t��N�
!������(G����K�u`�8KH�ēS׸2\�ϸ�Xs_��+K�M�1j��~j��<�@ir��M��<�;�ķ���HJ��)k5��� 	ףm��,�k0��/�R)\ JO�w��_�&ՒK� ���(�(�$�Ř/I��^$�� ���'���C��%{J(Z������h��+�E�;��v�ݱ�x,�}��
zl�}IC4`��'l�{Y�q2	�	�e�E�n�z����ė�J�F�(;Rw9C�4ҽ�>ϗ4	�P�.|LHU�7����A��1��%a�uEv���Zu���q��m�е����Ӏ�G.���q��Agޔ���cv�݄�o��X!�Y�H.RW�|H�	V��#1�}��?TE�)�娘�T��<4R]��'񈝾����w��o���ɕV�[�7@����@�S��|Q�q-�Xi��c�O�EP������槣I�>.3l��Џxl��l��!�4�D#�C�3�������˔��v"�� i�7=�����!73������0����6�b�b����N� �^򰝈�����Q$��Ķ�EA~� �#�_�L�����_={8,�Rp�: H2�NVb���n�}V��
��u���>vfה�_,�⛵�ԓ�[�\
(��m_K��̟���K#���P���C�/:�v9����,>�F�dN��w�����L��UxOw�=z֎�����S\��I�T�ǣ�E �F����3����c�&����׶|PL櫡�����W� �>^�������b��h��r>�s���ː&W[�&��Mĕ �~���dt�!��6ߘ�@�\/5�RЧ'Å ��P�B�J�����G�\�}��=�_�wi�Fj�g'������,=̨~~���C��9x��'|Ӵ��%���6�YL���7.|i闰�9��9g�ʡ�Ӵ�y�ݥ3��=H�*"��{�2N�Ze0A����Cr�ՆԘR$GT	":�����4���vcS���H�owM�;�#�z=*���V)���?��S!������c7��K�6Zl7� ��Q����x4o��0�,���T��ÊM�(uCD�w����!��F#�,�*�K���l�%��Ƃ��0��G9���2"0��v�$������2ƞ��U��hDX��L����b�s�j��6���'�?̎�|��KDo[F"�� r�,)�T�������H]qt�`8��B�I<��@`ܲ�S9����25M8�O��ܢGbb���y?��M��/\��\|:L�l��iо��(��:f{�]�-�g턑��C_j�};ŏC^!\����dC��z�@l2���uW�2b�H�S5�IwW}dJʱ^g���}�U�3�u�$)8���0�C�r���������b���Ҟ�:�_�P��|!ǀ��E,�����A��KZ���Y��g�y��l�0�^����Q���x!*\��J�0�	���17ʾc.�$����R����scg��F�mZ5�����lqrk����zV�����c^hY��s'��������4�á�b��ų���>]_dT�'�v3l��4=��r�ؐM-��C�+	7��f����+��L�ӞK��:�1y��A ��E�dz_H_��d��&,,�N��t�F��4R��V��ta�;]��Uˋ�(�)�TV��*j٬'7���9�/�@�k�#��O]ΛɘJVp�Ua����5惼Hq�F�}��<"�P�`�d��"�<Gj��0�BP�@���7U�k����؊��V�ib�)��1�[mhe�7)�|h��UJ��~��8M��"'�O�2q�!��*	W8��� �������CĈ�Q��9x�75t	��~^D�i~}����#9R����n�@9u2��P1*z��`⋅���i�����7�j#�t�*9D�T���#Il��o��H��j�g��i�*�oY�X	9�j]�Ն��Ba�Mz�	b��4�]��m��$4d*	i�r���������!$?:˚':�3[�3�����4R�+�zq*� �����k���=EC��<c�OŽ^�8�ZH<����?�F��ğ�w� F��������#���%3VV�c����qm)t��;b����T�`�ѻ~6��b�,�K��Mb��5S=��x����h�v����kzmQ� 1�a��T��2�y ds�j�hH���E��=�r#�(��6��aFM��&/j�aM�#1߷�hg��2�W��ԷZs��(�P��{[4��~���%���)����?f����	҆�C���eM�;�h���@	�����q�oU'����0��=UQ��-X$�|�.!^������'�s;����:�؇6!d6�p�X���t~��5?QϰcϿB�� �EL�dF���#U^4�yC����;��T^^v`�f/	�y�CWT�Ad늣���ߝ��h��Ă3��(�0�uk���G�Nn��@n$��gQ��|���7/�媓�iu�Qf��x�K(bIlz�-"�ȵ���͏���8�����㊷�'�WeÂ|�A���U����_���"v�v�>g������߅�a��Z�e���:�J���L!�8�bS	K��;�A%���R�j��w�Z���8s�R����������ӥ�c1ѱfz	��j~1����'��s`����u�j@��O��+�Zc���da'���M��^^�ޜ��g�~�'d>@��Т&]�}I�\��V]��'���o�X��_ܴZ���kBΎ:AUn\�y(�g2���Ab�&骠?�@�3e'�߮���щ�(B��֛<z�c�vF���S(��L#���k�j3��bs
�����R��Ü�g~`�H�Nu3�sF>RJFp��Nx���:����f���bZ�tnS��6�P3�'��X�����H�.�.n��n��+�����5��c*{��$�&�$����w�O�a��	�K&0aغǦ���Z����Z��؈HVU�1dF~����(���UǩG߼��댢��^P��"tbp�V��9�S�(�U-=�R�.���a�s�$�#�SB�H�:������;��IB��p�`jCy��\i�7uECŃ�RXQ+�V��g��S~A�Q�vq%8f���ep}�>;���x��L(���,�@}|&�ۆ��i7���xw?�T?��K@��iӓ�	
�$��pR��6j�����+��6���B�oR0c+CLc�P�-���X�&�u��ç"��_�?le����+��%�ڋ���]� m1��
|�k���b̭��Btu)�*\�y����`ls~����w� OiN��7qB���e���Gv���c��1��f���:�{S��O�����'�ha���s8��d=�:�Cb����wS�ǐ�et���L�z�M�;)�¤�F�Q4���	�?��MD����W\���66ho�@<�iI�z�.�W0�;�N&�L�"�D�<r��b).d�q�VJ=�Jdj	3A��/x@":_{WT��n�'��� 1����s�F�n���9{��A��ښL���5o����(��!�?:5�{削��i��?�x��a�5JC��&d[/Q@��+�hck3�I�+F��M�]�lX�a!8N@��m������<GN�IQ��+�Ia�i�_��[�J�0�͋í9p�� +�C�~��S tμlk�A�>�ӛ�M_���������i>[�;/�?ˋ<�bD�U�O!|���v�
� c��O<�y}��i�"9db���JO�z���Z��:g������+��X��O��HΝΒ�u�z� ��1���8�r��T�����:���5VY���]�Nb6��,�?��23�(`MMi���-p�I�0���w՜JMDè��7��0ʊ38��;o�#,3�D��LEy
���K'�z5��*p0
�[�� ���i���{��/�&���Fb�z�:��#s�mЂ��(�b�����M(�JD�����ud��f�R�,�-�Ն�uR8@h&�O�=���n.8V��tgG|�gb�<���A�D����7̗��bu�*�$����a[}#/���|m��V:���$zsC.5:В9��]�G|&
1~��ѭkc#�)b��>84B��F���G����S��9qjW���x	�1q�Ct�qi�&�A��'_�J���Z�Um�����Gx����QV���]zIQ6��d�v�i���h)�R��{ul��mxh�hX3 �X�nĈ3_��èg� �q��v���S]��N{���*��d���U�O�	^5a�#������P,=N(jՊD�zI]uٛ��B��`�p	[$Ǡ��E��F&���[P���2�j��m�
���.*Qf��̍i���B��*�%�t,���t�����/	�ެ���ַ�^��`
��I�b�_T��"��I��<������6w�N��9�i$�[��R�5��-�XB�\<?�uGluc�����~�ϻ�|9��<V"��}���,R�x_�ŕ�/4�.0T���9�]X�-����I�>���N��J!
ò�tϖ�DX�C��Z2����@�g.d�;��4�lt
�.E �%G%p����$�'�<o�"b !��
�����_#Zd�t`^Z�q���Z��/���顰2����A�9|���𣻆x3J��zp���Uf0�5��,%$��w��bc���DѬM�X	���Ǖ8�Vԧn!NJA"�A��Q@ڀL8��B)`�s�;�ʞ���]���H��ܰ�e.Jc�).���#�Χ�Bd~P��r�nbR���� �^1cN��a���fB��Ѫ(3GV�9V�)QmcE5mQ��Z�4�4,�}�U2���@խڱ�z�Y�V; @O2�U�`Ma�m*sXn�C�(��h�����(3��S:Ii�~��HjCZ��H�r�(������P|�F����畎UB7�Gwl�RV�c8���F��@D���I�V��$�}�r/���av�[T�:�FUk�U-L��s@�s͂T[g1��j���'�����o��p�6�3��|�k�,���׷��z�a��������r�u��ծ��o��Y�ʹ�98^�����fk.��ݴ��%|փ�r��Q]��T�L���ZXA�����������Lgc�?��I��Cú�d���e_��.��?�a��*�F9�yq=��eS��a� Bc�A[f5}8L���R�<kkEaa%$�p�-
���J��)ٟ�qrZP�m�10��'��q��A�U�F0?�Yo xj�Y���L,�m<��Ya#.\N\��dJ��J�x3���FM����$��뿦�s��u�Bv�t`͌oa��F�i�d����Yʿ��מz��P^�hEs:X���� fo����p/0Sa��NŚû�����uً�h6|P��Cj�a ^���1��= Y䔂�Wab�ű�RȊ*�Jf�����;B�o�D���Q�� N6���g�8�5n�)���a`�V� ��(<^G��MI���i0��NXl���LoD�0�+m�͉{���ᯉ�D���)b��h<1���ڴ_U#VРL�q|��T�,�p���b��D��xw�S|�����@4F��yn��*+)��t�+���ĺKW�2#�`��b��I����-ӕܗ+ c���^{z�%����"�\���Ɲv/������4��s����=th��������5�a�B�f�N��1������<�G#p^H�&UY�7z_2UL��T�G�.��,�p�u���ݳx��d�t�9x��"x�y�A)�Ԗ��,³�0��׊ۋs��ph�m��M&��p�-۪���v�s�(܍FxӺ �.z��}����]w�E�g@� �~���bZ�"O:swt�xi�����|���?��<*������Z����orY�8��fyQ�v��g�V?É�}�g���x�;#�������Q` `�fpPgf�;�3��L�%�4!s���oĎ� ����������̻��Nf��w�7��G�b�q�MдO��1�p�{V��!���,�x��q�����K'�g�aѺ���q|�hw[ף����J����濞r���Qd"6�ue,�,&���h,�+NPi#�����K�oW�.�'He��&ڙ�R�F���i����<��̀�b�D�G}c����ʹ�������jcFݯ9�Il̤������#/Y����ȥ�z���
�n����A5K��2@�,�FY�T�� �,h	�����tk��'@��Rt['{���t��d�N���`~����k��lW���h�J)�V�2���}	�ґ�S��惇g��������*e{a��F�tl՘Pk�h��"�B�%�G�UQ�D�P+I;��E^@�!"6�0X��i�V)�h�ۅc��1g���H˚��Ƣ�a/�D�-~�0v��_ �St_p���K�����-D��f�W��9Ƀ�Z�E]ɪj�j����Q	�H��b�7~�H�>����P�|y��S��`c���ͺP�ll�{��������IR���IH����?i��Y"��;��`3Nz5��۳�_��F>�v�Nz��~��y|���'� �$��'�cL[��ǹ�w�Co0��E���Fe5���d1��o�i�3-��*w��N����={q�������'��������3�3Qo�=5
q�:�9Opť�O��c�^�]�n>�(ER!���ؿ���9��M��јEmD=R�83]�u��-q7���ӻ��,���~�l�+�NO�N[�)���F�ݻ~V�VB�d�D����<ͻ,�m��tTo���Q��y{��rID�1$�v���֑�d���RcF�K�:�� E�-:�3�yj��vюxQ�����Jr&�O0Ul����9_��h�RZْ}��T�O`j`����<?�a�%.r��`o:�^������6A ����5%��X����;��T���?`;���$��`���֟��lN�X^'�8�g����T��}�umu�W�ۈ�9K6.��l	�Lݻ7���Q�w��$4��cv00��S�;|��nK��U累~�T�i��r7J�
�m�N�	2�.��ǌ��dGٍ��4@йHRg�p�~:�C���:����%��d����*(t4�XeM�_Lۡ��5�����E�6}hlP��d3�2��2�s
�N(@/�6j��L@//�i��!�����u�ذL���������߮���O�y��ԈnHk,p�[^'��y�}ۍ���'5���r���������:�vR�g�:`�?ll+9��C����@��<��(;��=���iq��M/"�������@fѾjD�?�$��R}����V�o��E��a���P�E�����D��'S�H�K���:MaC74�[`b}�v�����I�-����8�J�t�8!�:� �TٱM�j�e�j�/�O�k�Qx #sI_�|N��/�ŋ�J��I֐YK�����f�{�;G	?��w����U��4j�3��x����JiSI��CLw�"�T)���
�zHQ؛��m|$�I�&��2�K�Ǚ�$.�X<e�����^�11a�4:�Z�
b��
�����܊@��E�֗���l��P��S4*i���ᛲK5���f���"�8���Q �Qn���gh#��D�E�l�j���:�d	c�M��>֝l=�v�AYGuĂY�x>��'���Z+��K�,ka��?����3���ǘ�z5��iX�"Ɖ{��P�I�����խZ�"x ]J��Bv]��P�5+�s��CR�d�pv$v?��	��D^�v���iR�19��~+�o������2/������]��uCB��h���ۂ�(�R/������mC��uw}_.�IGk�zx��9������3�=��s)�5X;����'?4}(��/`.gcA����Uk؇"q��l���=]!Pk�h-<�Vnu�)�� G{�r$�ݵ_�KC���^��=�{��ɻ�B���Åo��^�C�#^7�x��HT���'+��@a'�f�z����"#��ـz2!�5E�f�!U!c��5�5��k`D	���2������F�]W��@���X����iɜk�Y�M])�Ê�; H�ߩ���cu/;,P�U1/\Q!B+�Y24���^�RZ�%T�n��8+uz6�_7N�՚^����
�:y+*��o�)�c��YB�֯��,�-ǌe�����v|�W��!L�#�	�NP�6�-�pG�FS���㣫<fB'��Q)N��U����/�q����i�刯���Y�|�t��y����k�v��8Ua��П)K��Ǧ/��,��+X�&t���)c:�����t
���3��#}���r<��b��.F5B�OA��B{n�,�@��&;��=�*z-�W_	ۙ��%�\�8��s�g{l����pvr����4
U+��u�_N�&�%���r�;oiX�a���3E��W@<Vj�m$��a��я��%|�"B ��1N8�MY�l��E%�8D�hLr�f�ƭ)d����J���h��*?�K>:7�ؙ�zz�Z��&���>E��AX&�7��[�c��\Cj奘@g~�V+��"�
q�e�Y��";l;�ՓXΣt���"�:���I-�ײ����Y��{5ߖr�|����	�V=�^���@<��h�P��@g�X�����vGޑ+w`鈦���69rѡ=&�z*^������S5��5Y�j�!X  'nh��z(�Ƹ�Q�U�oY��ZW�NYg_�.��*��g�e�o�Q/3�j�:���;��)!s�V��rh<�mמn�'���ӨB~y5��D;M�C'%���e&IQ��Sj�*�]^����{�.fp��^�+�*�ai������y/�^d�#Ѵ~!�蕁�揭0�)b�@������Xr��Tzgt*F3&�x`����Y)}��k��B�YT�p�����Pb���1�����T_+�7���a,�|k��i�v�y~q���:��K��;	���;��v�Dr�fE6»��mԝ�����
�Y
F�TSq[Um���<�Q���>�D1ʽ���@E>��)䞡�q/�w����=L�������R���#����(m��p"s��lԂ'&�o����/�,�!. �Nd�5:T��;��,�|뫦QR����ϒ��ق��X��]���=Ac�	'�2�G����'e䗼���j����d	�'a!g�fC9�u%��N�2z�^.��Ir@������vc2؍�-��j.�ZlCⴝ:�S�:nއ����}�U��7��:�B��l/���X�Ѵ�,�S��pW��0JlK��A͠��ԍ�ͭ%�z�Tj%Y 3�!;�9�8��-]�Z<3�['fn"�<�J<њ��{�C�
�e>T���5���1��۶$��#�ev!������d��
Y��ԗ$v��M�^J6R
tK�c�<���^!(@k�-��#�}����<%���'��ł�"v��r9��ܽ�	�?E�Y'zЅ��p� ��:V��Lx<�0� �N�����c��ס��H�W�褛�Lg$/�7�}d��}����>�g���X�,`E���<IK8G�AK�cw8#B�l���w��`��S(@�˪;�Ih���:Z��W���VZ�:���� |��bhqiKw��o�fԄY{�T��3��t��\�²%��P�	*׃:Z�5A͔#�|��!j���D֭:�(A��J�I�<�fTn���᪫���
*�DM�����gϫV�'���u)�����2[��nŸ��E]}0��K�"7E�� 4[���A�qJ���L��g�~G|_!뎡0"��<�
�e��s1`�SK�5ף3��68k�?�*�$�3��(&���
|�����n��;C����-��%�6�1�/N��o�P���Fb�cS'���8����BozH�,Bx�d�fc�a	4��K���dͼh������hG|��TU��-X��vsYa�&�Xg��S�q��=L'3ptX�A�J/7#���"�˷��q����|��N>v��UϮ!FoV��9m�ɶ���6����P:�#�n#Bg��_�0� ��oܣ&Q4\��«�������2�zNe�L��\֭_d���v�]�]O 6����cr������[���l�;8)R�Z�%����ϛQn!2|�B�U@����V�o��zQe99pt�Ё�ϕz�_y�H;��[�e{��<Xp�%�L2XKѸ��<��ԯsu��Š+u7�#6�8�i�D�y`��M�t�{�y
@�N	�D9��k�C��Vb\*��F�	M��#GT��7�&�&8g�%�S�!v��Z|%s^|�+���[ޚkWzi���W�����>3�ݽhW�DP���V��s?���aW�ź��'��EXv��fzs�Q���B7ؤ��
<�T��eص/V�B�	�t�_}Y��蛸�|�7p++�?Y?�ݼ[ci8�M���G�iV�`���#�T� R�Y��FdR�WC���<[�FB�tF-�_�����C�jH���1����Y�_��El_�0��R$:�2�	؝QpK�@ACJd�NG��6�C��Os��@�FX?xyPlp�>�CA���W��/��T�g��HٙȻ6]<M�q�2C+�"�yf��#��hu�8N�YC̢~n�H���y��o����ӿ���D�AB�`�aM5�Ю��!wF�;�1d�Ďm�#�Q�@�n����|1y��p0O.�7�3O���, @�>k��[	�HW}��XvB��ꄕ�4;AL��8�	�p�	o�9e�������a<5Vʟ4v�8��dx��'�#u	���G��v3W�:�"(��w
e~��?�_�ǄI�Q[�)K��=���'j'7�iE?�&��,�S�o��GPl�A��$���]��G�����@v������-V?�ߵ���s5�����X-0���lG&JgVSX:-�t d:p��h;��/���_�Q/����U��"J��."�Rz�Ok���[�
@+�1�3�%w�Il�T����F������2\Ԝ�9�?B���v�s?����H^˓3�u�K.���ܓB�p���.F+���Z��Ҧ(Gt�E����O�]ā�������-�Ǌ�$�	�E��{�Y�x'#�*~�Go�A�a�ǆn�M��O��-ֳV�5&��!c��Z����UPȌ�۽�������b،�;����;��K�*��+�����cf�AO���LkԒ�[����m�����)�!j�Y��b���������3��T3�e^3���S%p�:�#R�=t�H�v�h�ϣ���黥³���hLT���c�F������83�\���Q`����Ԛ��E�?�k?���bG�Z�G�R�
�L���[_�2�?���9����F�nj%!@���;p��"�t��9��䄠N*�
�[M	ך��޲�?i��]<�-�C�.�;%��zdK�k��p����_1�� z$�[x��F.��4�������h�,����96��'�!���a#r�c
�~;�-mGZƻ,���d虃F��}�gr������e���~�6/x�	��bt]i�ńZ˹�o��], ��^a�.yQ�I�?�񳿫)	��N	�ps��G�W'���"�FF����K��@9��沸|�$��&�<�'H�K�R5���}ffAn�z����?��*^��O=�3݂�v#�3aR�����K��F��:83`l�=��aSs����8C�����Nࠆt��{�}�	N�,�<%�n6���K��D�Kv�q@��f�����uJ3	E������	�2��!��H�)����]���d\��r7yw��7�ʪ��0��4>-�2�or5�0y'���vٚHz�ط����5�b�B"c�/��8{4H?!-���݄
!�-�8�9�����(<��RV8zs�7ʞ[�B&��W���Ƶ���z���i�5�t;qa�L)�O���H��n]R��E�k����h?����4d���F5n��vdQ�j����n�����T��Z�r�X8��T���1V�$3Ze.������Rƨ�{��B�-~�s���4�5�K�Y�h�	���Q�`v$;%��d0������-L}1/�vG$�{BX(ǌ,�|�:�0<��0Fԛu!�R�'�X91��}�7��Wh�;�� o�Ȫ��=ʶ�ͣǪK=�(� ����RL����f�l$�"�n�<��Q6�a���yO>��X��t`Ôj�x�c�����@���-y~����'�{Ip��S����M{(��E{�� �t;J�F�;�.����$��q�V�pë�������^��g�{b<
����@�^��R
�)�z�?��>���I�&U�x�
O��ηK�='�މJ�0x�#H�@���>~7G��K�Ĳ���/����*�B1��ƗA�E�PVq��ԓI�{�C�+'�d�qz��c�����N�����ќk�%F��Yߗ'
'��{o�+&sR�ݪNQk����jQt�k'Lm�\6���4Q]1����}�s\9�:����ÕN�����,�� �>~�@=ZM�9��HMzv'i�w,Ft��,n�;Q΋����Q�=�O��&��`��� a�$cU�C[�M�l�y��˥s��<�[>.��d>`0:܏�m�h$�v�h��R}�d������b������)��V���4!zS<,���z��Ϡ�3�Uq�b:`"~��&f}���A���<+��L>a�e��Rmx��KH��7z�,�#a�yW^�`��%|�r����9�NG�T65�@�@����n����()�࡬'�3$K���g�v�餟�ӑ�cc|qq6����t��<��a�'���� B�`��7g��T�O�f5���~��`f{N����>[eۆ�'x*����<"����aF�����Z��w����
�\�m�<[��=�{�k��x�8ڦ`�tc��-oAL��^=;E����kCً�,* �ƴ�?g��6��(��~�#�z�t���]4�TQP�=u�+c��z ��k��,r���=ƅ�qPhÄ�C�&� ��LZ��­�bûm7�t�-�~�uQ(�P���|fT�8����T��#��V��=�]�<�;� �$�4�:`���c�������;��j([����*�u��^�eS�]�{I���&*`�)qSM���/L=щ�*�ܻJT�-��)����K�b���M=�����9�
\�_F`�R�FW�t�7��{f�r������ɱ8��C!~h��v�ˣ�*�*d�I��(��?�y�hvpH�������������fhǛ�zj�M���ܞ��Rz�Q<vQ�byS
�F+�����e�rM�VV����l�"�o���a�3�d�Ȟ��zT䛾���E[:�E�%�f��?���h�"�Z8���B�3sa���1��R]����t�뽳b6��?:�K�&'���ql޿&p�,0��_t���cI tB��)L���@gy��53���jj���c`Yø��d)��:����y$l�T�T�p"�^�=p&�&B1�P��C�]E����/��D��m�^��~��:wc����fq�[K+�%5`�b�[2�e�#��La�t���>F	_���k%5u��E>��hN@�GW�_ܻ���ʓ�l.�������?~�����ML0���)����K�&�UW����0��-���M͗"ir���aWf]�\�'[hP��ɱ���)�;��/�F �2~TF��ͶX��e��M"3?�����m��[`�'5�b�5�	
*��/��e��T�h�V \KYP�{�%&с�h��B��6e�b��
1v�D��wJw�#?&�r�G̉�M���� ��p��R8�)�zo��-rlŋ���Xp_l�wԶ|c#��>4�k�Y��qR�d��s���nxAr��d#��|�ʹt��%��0R�.8ق"H %F��Z��6��Z�����Yߨk�ȑ�Kk`i�.Z6R�����q6�kR����Ϝ�\bl���J�V`"�� ����5/�aU��?=م�4�@��
:x��gDGLu�Pp/��}3x�Thr�9N��;x��"zt$s���Λ�D<QmKz���%�fa�K@��{J�Q�B8�gq	�w�9�䙦��.U���l�����a�a�Hr�I�g� Ya��1�������%�fI�yY[�?�7���M�a��ܕц��JI�b��,-��yFv�F�DZo��pC�:8�1�NF9�!*�dX�#�UQ`�Y ���ZV�J>�&ǐsHU5%�(o��C�ZB@tJ"{��IȮ�¡���֫l�'�Gb#�Uv[6Js�Oʵ� ��]{�<�O�-5Y�Hdʨ��d�q76��g�v���t�ѦD��(Q���ǺA(�!�v,���B�mj<���yԦ�x�5E�P�id���xgX$ �f��&j3��RU#�7���[���V��{��J�*�{lx7�ci��Jx�C8C�3�H�D�0�+�'�:�As{_����+��T�G-8��!c�u(7��޽[��Oվۺ�l�YA����m�R�:3��?C��h�7�c�3r��Wu�|��
�Ղ(��� Zi���u���\�"�����@��%��7T��y�Y�)J�����z3�1���>��?O,r���l'mqo�<�dUz�fx`�0e�]��t�6��H�B��{T�`�,+p^G����a�x*�c���T	�b��e`�W�J��T�xU�Ӥg��Y(d��>���F� Q:�r�2,Gk(�cb~RY/��vB�R���\{�J�Tdkѫ�_R�I�'^f��1ED�1������ ��xdL^��"�ׄ@�К�/J��w)�<��
��O�e�6�Tg1�5�,�:C=E��=���@9"-�-2� i�2R� G|<3Ó==�+����h���dqɋ�ɞ�~�Mu�?��դ3ћ��f����*�?�
�ʢ*J�J}.�_I�r��9���z}��'׺�[��n��y#��Y9JY7c���V�|� ���ش��ŵ*t�87�M=Yn����VW�O�i���~ܝ��nXsx��E���;ظEX_2��Z߆d���:�/�����d�'�ÄᏉ����$<��ݓbq���]�.��҅FO�f�,8MO�g�M��������*�}@,���9U�rM� ��=��"}��l���3��~��!蛡�䖴���\�|��[��e�aa  xjyu�#�,f�e��Dch3����9n�w�����P��H�@g����rV�-[�Ū�ЋF�.]b�N���+��{��������R��;�H8�x����=�����S�������tmG���g��A���A��Yn/>��by�J-�A�2���8�DQ��x�/�_-�� 6�U��%�R����vH�G�f��1�S�R�!v��vŻR�����h���<�)��"�n]��"��,d9�{�af�>`�U�~# ��&`xq�e��,@����7a๿!5H-4�X!VL�j$K�?t̨t���ڋ_LVm{�qq�,�wil��C	ӡ���ƭ�4�J�O��-A���./�I<ˉ�굼�g�ǁE�+� 0���Q���C�|Z*f�e��?�j��۵d��,Y�<��Sb1g,O̝J&�� 4����r����@ٙDi�aYId_j�l���6�!]�)3�N;q�W�>7]z���@;T������jnwA���#%WX� �nr�,*�v��eR�iL�B?!��Eإ�U�3�`DR�zWVo��*����)�`*�[8�GX�'��o���'� ���rN3�c~�A'n�}�Q��l�k�AuC+�D�L�����	�0�k�eb�ty���8�����Z�5b��`�b4��"�@gL��(p���'H�Y-��X����kB7K���ك����_���\�`S�1,�x<�B�M�t	a��WZ�936��s��	4�Xɦ?���YRL�d-��f��筹�)�?�i�檕TX��";��x�|�9� İV ��6M3�aO����ʥ�_\��LRHUU�
ds�������V	k2�Β~�qr�M+dr��헸M�T� ��F��~MBd��M��2�enh^�q@�f2ל��z��l ��*���68I�,�a/"=�l'l��p����L):"7��r�7��[�"�(e!Nǔ����g{2=|�u~�:z!�L������g_���m���^��{}�� j�0[��HҜn������Rߑ�G�a����XR�g�S��7�a��ެ˰��q�	-9�՘_�ձl�Q�֔^k� -N�}�a�q�i4c���;�2��:�-��33�Gezҿ�k1I�m�K�Aߡ�mQhR-��-<��@H��!�&lү	�����XR9����n��w�%�R��Ђ��PS�������Q#
+}��ES�91��q}�8�6������/g���"nh#��z�,̰'E�ȶO�n�W��:@�~u��]��T.�.8kƯ����j/<��B»�n���si5b퉟0
��;�8�m캁jgX|rTx$�նCΞp�\)�{c���T�P`䤋���S�஄����I����;�i��-5SX�g쬴
�����z�׆S]����Y�����X���#�����o�n�[c�
,(/R�Z�+����S��p:�Y
L</]w��H�;.5�_o
�#��A٣�@�H��Z<I��J߀���$���:�C�sr��V	 %!b9��@��\���#���g�˦Rg6��]�) ,.�!x�α�M�b_�fWʆ���i�(�6;���	�<�)|t���p��V��Sox���ؾ%~�r�qw���@��p�O�]<��t�Ou� .��]kk�C�۩|W������@&��T��U��>q�WcZ��O���#K+��R 7{�S`�;-�RM�@�Q��~C��x��ڬ�@]j��F���˺V��!�uڱ�4K�����ad���Ԧ����GA���"�ދU\�޽�N��ᛛۢV �G��(5ˤ>��$�x ���H9�%m��yn��l�� %�٦��!���8�F5휑.�Q�'לo+���˖���8�Xd��,��˸���o�8v�Pc:d܃��0�#=�P,�i�w�< ����FO���N�(v)|�K��:�L��0�^l}���_Ǿ'�r@�]�4����|,١ʭ�<�����	�d�\���6r�#.�R'�Q�pk(_ 0�gb�]�/sf�^H��#��	�A[��e�<?+K�^0u�lS���\��ۡډ���do\��#S���Cc���fsa�}dQ͚����*TÀ��R'���=�e�&ѠB�����x�x���u+���i�ӟԄ���@.qN�i��VL�F��y��G��񹒵�����a�+��"Y�
�E��IÑ�L�N=/����鲋�r{,�*�}J�/Y�Fj��8f�� ��� �b�֝�Ęf��gZ���ɯ[�^��`����N���J����n�x���E���%�Z�aA������x���"����;���l�]k&߰pYڃH�I|WY��Wa��9�;����@h������'�9^IP�˱_�^�NC��v�çTm���vvf�W	5U�ߨcB6/&����-�q�ϧҁ�� ���筯I���-r�wAw0��:·��
LCAr�8X(���:Vl��Fzi��)��Y�uؑ{���4�Tdg��M�I:�ZH���B'�,:ץQ0)r�A��7!�R7J����^i����I�1We�ϋ�^��Y]��gGx��]5��A��I٘�i+��I�`�H�M�F~)�"9�=��>�W�z���d����^�A�Z��w�t�!_��=��k���f-��kߨ�(�Z�����K�����ߌ��韢���^qW<n�:�d��mt��h�)��z�,Hb� �0T>�MH�v��9�U�����¬*��A�����SJ߸6���$�S_�$���
���Û��ӳ��%�ꋚ�cv�'+U�nū�O^��*ؐ^�{��e��t.�p9�z�oL�F���PN��x�����@E�v���o�O��1�n*�";��L����ǒ��v��"M:|^d�
3���T@T��ZI	���qX�����bT9QQ��ͥ����7j�v�{*k!�KYbd��*b���g�%�ɸ1� }�Ĝ��y����,#�t ��v��{=���x|5Z(�`�I7�`q7�$V�-J�d��Lq72�܏��r�G��G���5i�z�T��h_7T�+�m�����<�3��'B���L`��uS!��R�5e�[a~��]:񃢊���OHK�wg��y�=���4|�����S)N��K����$'|��ej����z����buU��Я���p�cY�Ԩ���
|( ���5++�ۙ�߅�}���k�?޻#��1$�6�]�@�9j{k�Lvs"���=b��n,	ԚF�F˚V�@�gΘ���ݵ�h1/%:�㙚�g�z�]�c�yi��H9Gu�k�z�󜋡�՞��\0��:8���:�g��N4�y��)�o��]B/��5���m0X���.��-���5���6ya��m���D�ke޵[>��*p��c=��
��ց��O�	l}p_#6��@�&]S��&�m�U����U��@�|\
#_�sN^�!��I��]�@1��Z��vV9�]{b��ƨ�b�����#zU#��rg�X�h��<]��5����ڼ�f˿�#_m�d�0��?i2)��c��x����rE��- �E��yO����|Q��`:^��$haO�5��9?�}�-D�#�)�OH�ׯ����R�寭&�|�;"�'�{��ڦ��VW������Ғ����o��Qx��,�KHm�?����t�|< �D�����xs�w_�,/����{�����з�x�rB/�Q�1�5�\��3�����C�#��m��A&�-�E˻�S�&�s�+q�<����^gh��J�G�b[��['�A��&'�{�^j�y����Ԭ����ݏ��`Ć��d������9�ܵ�0�}νT�F�� �����Z�~ܦ��M��d��#j�ek��\vV�?�G��Q�Xͷ}2
��%`[�ׇ&U�G�"li7`љz�AN�P�~�W`'��麒�g%�2S�=�S5c_p��� 
��Ui�soU�6�{����'�+&�� ��ճ�BZ�f�B�|�A��߯�W����|����=����=r�m��,���'eA.���F��E�5�͹�O	tB���r��M8T(s�P��`a�t���NO'IӇ=H��}���a7V��e�t��q��AR*�h�)�eo7h$7@f�X�m�K�'�Zlo�H�uvzko��i'�{�X�#�}�+*���*�Պ]O����9�h�K��>�,r�ل�̲;|wK��M���c����2�t2idq��^xdN�LF�F�`�g���Y7
zbʬk&��gl^R��{z�iX��t���ڃ�}3`qs6t��*�����b��o��:�š��)6���X�k���,(�u$8�)-x��Hfu���/�Y�q��8�=��
�*�l�*y��t�U�6�� 3x|�^k�:R.1B6s�u4.9�/CXa�*���֗�Z����a��bA9kc��|����V�<8��ѱTB��HBX�T��AD�����:�8�Jʊ�����VL�%d��)��g��4l���?S���$��p��w�v��~�u�X��k��u��d����F�F�h����Q$�"xl;�G�7����$-O�Av[]wIF��c�XF�u��x���sy�ɘFI��y� ��	��j)����ɳWh�g�G���9Br{P髦߫���v�;j�:�Hsv�Q,��Oq3b������ZQn��a/���T�������� ͼ��G�Q�S��X$�Ɉ;e��~��>'
DCB���nQ|����'�~��b�*B5Ѹ.<§5@�\�10���S&#������`%ļ���AE`l7O��W>�chfU./x�utS'�����k�!��W��w*����Z@��E�E�T~��>�����:�7����qc�@?��Y.���F�||�����ʹ\�v�ܰ傱�-�H%��b��� T�EnªKキ?�ѷS
Nca<�jt�p����~MP��0а���qIc�#���b�<�������_d�#h�~���b=��Y4[qdu���b>���C����U5G��������tQM8�i��X�^�oٔ+��1 8��6nWo=��C�����0�'#'�u]�=s����k����|��(Y̤�+:3اF���J�!��O
MҀ�ܵA}Or��4��T�v��s�8�)��bPrc+�B����Qn� �x�l/ʳ�T�0�b|Ҝ�P��#�~*N�̨�8�G���m���G�.�,	�0S4x�eVg�f����|JЏ����6m�aexѨ�1e�߅��x����O{���ξ_}-�[6D�+P����E�����[�y?�I�3~�狋t3�J*���c��'S9�ly�I�8UP���1i�΍1vC_0����������H���],�c�ޡ
N>��rG;Sd����o��7��=�D?�%��*�2�.��u	ߕL�x6O�cmK.�k��zέ���_�`��p7t�+f���y�y���U{&�e���x�+�2E;�J�+gsG0�2�t��%;q���;�K�,W[�P�p�����?��Y@��uZ�TJ��:K�{�� �#�3�I�:�v	a�N�#v�$��6��Ͱ�"�|�GU\ԢC?W�����k�ҜέɿnR���С��ߗ����2�
��enx|�4��
���tAp7VW���s#\�����&<1��re�����vH�{l�K,�����'��,�N��P$���l�ٰ'�2�0ܾ���&��}�v-��U�u�������%K��P�Nu0��ȯ�� njܗ���wyV��i���_G�2��PMa���c�%;����|r@��).�ա�kq�"�N�C���Ր��'���A��
� ���������8B	)A�H��om�������3��`�YΧ�c���ac}8��Q[��g�����? p�����8NC�,<��=���$��R���M-1VgƵ)
2G��������jC���*^�]�e������������X��4�qs�ZA�������O���q������
�`���J��Cc�s�"{P��D�x� L��I"���"�48�sB{�����Sn٢�o�A���:�
Y�%q��V1Q�m�TR6̡��d���F�%�q̙��ST�g��Z*��N-X�U��;K�ב���U+� �g�E�dG��5��]ǁ��C�Z�罒�*c_�J���H�sq��+�-���x��Ϯ�y���+]5QmsY�[��4L�WC��R~`�n
�a�7�΅d����.��K�h�N�l���'�s������N_�������V;!P5�*��~JKTg�j���!@��8�{�!����5�ʗ�t��wQ�P�5��Wՠ�����/�W2+��T��gl�l����7��0�Ja>05Hf���]u��̶t��P!�Ѩ�j�wC,�`���M���^�,��7ۗ����b�o�����|�%IXt��ir��,~R|kJ��1���0��X��ƶ��]L���6�7�o����.w��T�e"�X�8�A�n�@WQǆ���CO	�lש�hZq)՚J>���T*G [��hO�V����/��E\��݇��-�eݰ�M2↼v֗��;}��s��{c��H%W�,�'�+N����g*�s-����	��o���@���b=^PW��Fc��vTHurd~6��ɉ_��<3f8�*Oz�1XG�3~�.��H��Hxq�t�~@yU�`�;_�v�����<gV�Ui1�I�K���H��>سp��4�/���!'HOq��B�~�r�V/�r�P�6v�5w��:��/ ���?�ޢ�V�11�4
��f��b;�U5�.?,P�
J��_���.���:���h�+��B#j�1�
�єB���1P�� ���LP�BDt��˿���@���}����|�0�\�i��5�����og�v}~1X�":�/7.m78	7}��.�����x�~�]�UG�^b�q��iS�YS�|i�M�K'��9�{��V	K3#�|�H��Qd��]5����2to���wN�������F����<��~K]*�2ظ���z��FU����v��ߍ�s�g������q��;�,`M�`:Ǩ/$WN�Z��L_Փ�i|e�ׇ	�Bq`�vK�z�{�z����X 2:n�זz�w��E�d��~�<���3�\�e��*#�uAT
�V��O�AD�bº�i=�y��i�7��6@���p�Cj���s?��[��,ywS�H/���]���I�[?|_n�(�R��[X�;��^m�h�p䞑9`�Oaz���+�nS�>�rj�tր�fw ���5|���Q.�]�I�Y�����S��f��n����|0 K~+P-	m���m$d({�i�i��D��$��Y#ަ�X@��Um �\C ��Rh�I��n.X��(tYd[��ڻ�����/���L�U�ʍ�(�Hes�b���� ��;������Ma�u��|4�0��=h�����+� �J��,�-����xfKK�WƹhZ�!Ǹ;����(�7��5B]M�%����zrS�bU���{�JI}�Ω���= �R>�4�o���_�՟INX֝�	�=+���A{\���LX����a�%�]6�б1��3Hن��o����ȧ"���W���'�1��F��)\B��Ng�.w��w(��0z���ލ�e?�����?�~U�R��'oϼ_��{�&[�Xu�� Š��֋���'~e��ˊ�'�{ס���n1h��9Uxl�T� ���.bu'� Mh����v ,%:D@G�ۅj��ty��������F�����ڟ�{k�UXx#t'c-�{͑?/a\�fC��3|��|t�X�>%��}5���ܻ�ۉ+Lac�Xfma��59tg��� ��������?u���N��>#ز�Wݓ�B��ߚ�}ޱƳ��q�4�V���7�\	1k�����V8�kH�t?ElcU��T��뤔y��R�)3������Y�{t-�e6D�<U�m
���z��R@6�[%-����b^�u���)��<`&t�r�&=F���[:T*��s:��N�OAѳ��/��'u�T�����+Np+J�ۦ��a�_�L�ه�J0�s���-�������i5R�_`~�c�ݫ��;y�L'�πZL�#���>Vk[�p�3}�똶�����H��L������'�ӛl����T�O5�{������:,�Q�X���tJX���79td�g�S�.�,�W�}�`��0`����P�q+P������m�D��D�Py�+'ɝ�zX��H�Q�Κ���K�}�d�Y�P���)v���ޯR��5�6������y��"D�Y��f[}�ן�/��w0�X	� �>�(�>�T�N����|����q�|{^sX!7)�g�F�)@LXpT4�AP���c��NQ�WA9<���M�&IVR�5�?��Q�	c[RFL">ؐ�f�!i��jZ������4� Am��OB�xV��j�d�����vv�_�0�l�?j2c��D-���:�9&��F��g�#����-�41N�=�-��e��@��uȏ������J& c����ڍ��Yw3��	�ë��Q��_5��o
TMJ<���C^��I�'�KN������K���g�}hU�)���D�>B]i-;E��<���q�=$��� 8V��!��dTP��9s[�!��u�Ζ�Ң�4��ȩՆT,*��~���W���~���S�!�[�`7ύ���oBMu��#ё�����p�ˍ@��狅u��duH$S�0N�,�!eg��:'�)9���z�ptB��6����y!��2n�*R�C{3<���LW� j^�"M�I@����t#�|�dx!���Bcτ��/ul/q�:����[	b�J,HH6b"6hn�9)�lR��iN����̝'�fZh�6�Y`���Wu/����RVը�/`�q%h �=��Ѽ�{�X˹��2ī66��=���s��(�����q�ɸq��Kͳ�	���9x��V�0bO�.�atA=x�oY�1���~��s�g=�i3�)�:W�'��Rq����� a���ٜ�ȯ/��&��?P�W���N�οO����F���]���l�����u�\M�F,rw���VN{j�5��x�ȇ�H�T�;x5z�����MX�����ADWX�\�Ӌ�����罁���H(��y ���N'E�����Bm��G���xEtx$��6�NA�����`�Jk�@移�<Άk���In�+a���sRR�"�<5����o�<�5e�YLП{�7^� d����B��v7��\9]&;���-M?9$�aa'�r���1<u�A����H�ڱ|���Q�����,GY���Q$�������1��yӷ�^�F�����BŭN��؝�
��3��P`�Yi�~�Ǘ6/%��f5m�����f��yJ��-��`��ȉ�6�V���Қ0Ԯ}0�T�4����e�I��;�x(����7��Wīl��ڱ�V�P�v�xL�9��R�Y	�t*�Z1���w_l����M�<�J:�����lr���}���V�0'����s �|g��H�H#�1.0��:p�!��#v���FQ+����I���0�ҽ���i5�Ϊ�0�Gj&O�����3�?ԩ�r�b������0�Yi���]t�hX�1��KG}�Z�QV(����')e8�U�s��~��7ֳD��#g�b���QJs�.6{+��n	3���%���B�H�(�wq��X�������`KSƋC�_�z�"�X�m�]Sg�,G�{���b��'��>��ۥy�"!��8��V�mA-�:�@G-v�>f�ms����G6'�(W{bSՐ���n���	z�%*���p�=ݷ�4ޚ�sSH|ZO��X%��@��ڧ3��G�P�"��lP�DI��|�$n͇�Ƭ�� �;L{��Hնo��1eY�fJk�kM�o	�$gU~�I������D�,�-^�y��;%��d���d���t���L�T�_��Zxͼ�$R�J�8��>�ě�=k<�K����`�|T���M�k����I���\ �)��7E}��b�O��vޏ�T���w����?���ޅZ}�ɟ�\�����!�r�@G�Sf.[��̟Gw��74���p�"|������	����_n ���B��/]D�ֹ>��)k���7�U��֕bw%}p�\í�U�v�w���_6��d��+���d)�묭)=cvU5F�		�&��y�/;�^�:"���-�ŜR�=����~�C���fI�H�4�s��_��ڤ 2��"Q�>��)�����2#,�Y�,�h�����V�E�~9����G��(#�_�Cs���Dd0���D�
��zP>q�-��7�KG�I�b�^TzVBt$����I�s���Z�]n��������0w� 8��T�7񴤟J�P�I���V;)�8FXJz�mY�J��jbȵ?�I�pg�WR6��1���ɽ6�-2�9�C0�|Q�:�T@��SO���N���(��h���b*JDX��٣&���:!�"[�v�>o|c�ͫ���w.vx���8䟡�)\6�Ie�b���DV�Ȃ�&@ʽn��D�N�N��Sun��Ι�(M�dV����2���X7A	Z�}�W�?���Lx���Wēho��O����I)X�u�.E�$����8�S��-��a�z��Hz�
�*�A�J���?�[@aݫ�y!RO���5��?3W% �%��hI��wme�!w"�ēM��,�cR��_*���4s�X��� ����5�f��7������`` �͹(_�[F<璝����*�J	���(*R���K=�խqt!��Ͳ���� Ȳ�B<���E�&!!��$`{�!�K^y�a��;U��&2�[6J��]������n��,>���Ԇ��H���&<��kw{J��):=���b��i��c�,�qd$���h��J�xH�3薏m��*Yv.��8;Y���})�d��x9�NT$��n>Ua��}� �3��Q���`���n�HDo<�~�<�$����+��6��E�!�>� .-�mMTŗ��^�i'{K�sY�P뮅*; �Q�����#O�����[3�
R_J$|r VP�X�{ӵ�МR�P:���$i���11g�����|��V-|j!E��
\���EF<2��+�&d|cѠ����u��&׏�[�4AY�3]:�B�E��`�nhy���5IȾ����̈�R��qg�.�Y�Z�ޑJ2&(�:Y+RXpKb���k��8�k(.����(X2�	��E�þ�T���Y��	�6��Y�׿8֕��G�W'�>�E�Tx����t�x�T�j��~d��>�.F-EH��>QKa�z�o9�L�.�gR�<�����HF ��S��5�ϼ�8cY}?�~�X�&� ��<���*y���}���Rv�#�ǯ��]�3����Ӽ�4#�TT�D�J(^�eg�}�[0������n��ܥc-z��;m�ve�#��2�y�ȮAo�l:��XL*(��jڕP�w��s�p�O��v|�g�0�ݤc�T�N��{%��<F�����14��Z����%AB9��E�AA���j��bw8�z� H��}� ��>���*Յ�Re�ػ�C�ӗ�yc�̙MA��@���X`�V�g�(<�� ���,�u�(Ǽ���4e�2��|ط[ ѦԼ�[���1	)nK\��v�ܓd2ݫ2�Y��x�~�@��CS;��b�!q�Bԇ��t�+^�&Q�\
j���ǩ��=�L+wx�������dY��`C�L{i�&�Q�>c����]��IăT�|�������r�]6`����}��V�Y\/�Qh�I���pa���/��o�Y�zw_k�eu��zz�%Ɨ�2������;c�Ng��l���ó��R���2 �S�T�GK��̅w����ι�\2�T�j�4l�ih�YA�U��uiJ��f��Z��9f�W:�s^�w�:��_�&��Y�$�5�;X�g�<5 H�����ޅe-�U*�g�k�p���u���:F�P,4Rq�@}2�V�p�$�8� ���{���XJ!���g8X!�%�TZju�\����<#G�Ucg��[V%�s��kP)T����(�!�nڻ0W���2QHr�s�<.x�ځx���}���9���1���'����D<���0r�}2	��?�.P��C�����@%8�Fv�0������X��~e(�f�"�@z�����|�-".}�_j!�
 8�f��o��e|�9�u~$�cW�����7���h�JX�����T\���3Q@��)H��B�x��醨�@��<�����)��wrm]g��M�-��V��� ٳt�s!U��nCk֓qĭ8��9�������#G�05�#G��?�U��s��oF�h.��0f��e	}������mWP�����{����pOO���H3���[p���{&q��@Pa�<9������Y��
���l[i
:;��ē�>�_�,��=/[�
G�25�o?:��K����G><5x@s�c��JA}wѾ�����QQ�TC��j�~`C�|�^6 �o����E��6�{��Z!;>Ǜ1Á~����nX�svcɺ�iPu�����	h�!�4�{�2�N��i�3�C'0X�8h�&��c��#���O�s.��e����l���݀kp+�xKL���v�j�Cu���/��mE��ǃ�����ʄwU{w��^N$��Ž�\[7"��V-��e���ӯ�#��-,Uk�FK
�b[T�'\�U���ݝȟ�%ă�������s��G�>���H�����/\Q=��	-��<g�m��!�T0$�I�ћA��E�+K�����EE����&����F�|D�}�RXa	�n�,=sA!�=	n�Q�`����k�iw34�|�bX*��m��t�# �t�)�[�#�Z���m�u������'��"BO�Ve�3���X-[����ɺ�e.mo*u/,�b�lD�-/_ ZU�ʘ���l�z����^?�U�x@��ߑ#K���ګ��c\r�.�� ��$#��&�P�W��~8$�q5Y��v��CXbT8����	fo�9�ө�+���� ^�cS��F�}�w�.h����{H#8d�g�.Y�slr
�T��td0���N:h��z���?:lĪs�m�!�i�ݗ�L�}0���F��b�Ve�I���Y���Z���μ.�%�;e�ZEX�6o��v#�̻���v}Wrq��]������;��D8���U �_G���k���&[�׵�I���1�o��g���N�4�q��7�ȭ0TYr-��F�Y����#%�"UI���#N1~ei�9��6�ڹb�,|r�/�,YFr_��;��k�t)���Ԅ�X(��`���䪐SE;V���U�L���5�?6]�)����Q���ɢ:��$u;bd�p����>]�#���*}'"��Vp���Y��2�_B�?�2�W�'��*�JN�H">�<!�����oԷj����Iu��)����0�z����<��ݰ� �BpkJ�H<r�*����GR�D�~i�b��� Kvm�憹�C|�i�Z���gE)	-���J���F`�<�ʈ�x�m���Ev���|(\��k�<���j��a�d��$�>�jN�2��������� �Y�˦B�	̀t��J`q�(��E�[�Q;�elYhb)O6��ټq/�@�}�ʏ&��s�H�or�7�y^A{}��^gyt*1��`�?	��������jFF��%&]�)�)�/Za/~��f+f��7N��;p
�7p���m]]lи���[���٩q5����*7�^c.tW��״ipU#����Qf��k�jp4����Ѩ^�|�x���ޅR��c�xO��ǏB�N-��{��	7>�T��;��� �����]��"X����h�ʺMa�.�*��I�}�H��g��ǂ����]���e��5G�{��3pzQ���m�Nt�1)�G����+��Q��d�7��gIa�ه.���{��}(���S��>E]n��	|��僈S)�ɭ��8s8Ɗ��JX���.�Bu�uU�r%�d'��ޤ�M�܎d���dAB\杰{S��w�p't�8��ʃ�5�<�����,W>�ޞ4���OLiDg�t�z��Q�@cP���,ҦU�EP�]�g+ά�k
`�=5ċ6�Ra�w�E��P�i�hy e>K�(�
�$�b��	�S)�v'�5���}���r+�4���m$��Ũ��w䷁�L.�x��B�<f����RJ��4�s�t�C?���`�*d�)5i�tN3����_�}yo*���i:����%�4�x{a��2 S�ь�f��?�h1�ϳ��!�#��$c��E�b�%�L�gJ1�Z���+��뗪��=�ūQ�e��)���D�J�
�@CE���7�_ƨqujG��U%���p3 q��F�6+���V��8կ�7Zk�-;��!��a�	�TǞ�mC�3'�w��Q��Oo�=��r�Q ����4Cxh��?��B��) D(PΨZ�6CB~^����r:>p�.�������o|���ap2d~�$�e4�X��Eu�C�?d�З�����cm~��%-h�G�}�2Ks�auω@1�d%0[	
�0����D�bM������'8,������d������TF"�Pt���Mh����,4�A&��q| ����p{H���k������e�!8�'��UF�(b��L�.
)��z�i�x�7{�(��
=02�SBddp���OVK���~��k��`4(h���AUs�$h�%���d)Rn�PŶ�B��WŚa�:_�\�b���3����K������":�-��~[h�:OsUQ-S�����4	���~�.�	'Dd
,�^�\�n�7�4��W�w��@q/SZ��rY�}�C��I�l\�N�����,� aR��7�<
�6"W�����������3�:&$�O�>=_>�;J�wV;$p\��ؐDݢX�1n�\H�;#�n՗�>��b���{֕F�N~A�BBU(I��b���X&�p9�t�W�3��p� �7[������d����%b(�!�8���"�}�:p��[�{������9�9M�������:��"���ֿ)�/�wM^�&�!���|�f�ݦ�p�\W��7xY�A�_��e�:nmu�}�c-/�~�g���2��`�xL-�z����i��E���V��������.�'}�:ilǈ���t�<��g@�O� �k�e�?
��rU1]��RB�6*�ͦ3��GɆu#���e{��������*�*�9Y�c15�nMc	ɍeg��2�Rֽ�5�t���x_<Byz��ukj�����ӑ�{�X�ڄ�\���ly��.i������v�8��3Ufi���G`�Yʹ�.W���E�צB���$����ߟU�(�y�F&�DGI�O��5�l���WG����;k��'�bgÎ��W�x��ג��?�=�"�6�"�����8�����Ʋ?}���Z�g�s�/R��c���'��u���%�C�,��7��\"�gX��z�C��y�\� �c��E	l����vׇ���D��)L2�Z�.�'j���+)��]nU�V5��RQ|Z����+a��QBz؋��4���5�a䣘���f~D��M���":^���	m�){����k���\��8A���Ov��Un��d���[񸬨$ND�h����.���q[RTi�?�v5�P��E���k����1����St��.���C���Q~�RcPl��^@l�쐻d+����p��n�ⱚӍ����@�SWu�>��{홞l%�}���kQ���' �Q�@d�&4cI���5(������|̍�EZv�d��#u�j�o��cn�������:@'��`��Z h���U�c���FN&=�E<�p�b#��NV)��p1֏���ۧ��N��p�����>� ��g��e��kK4q��䍈��l�y�fz�S���K;���r��8�)�������HK��}O؋���I;�O��
U�O�Ee��= �TNFW����E���О���t�@y���=.g��X�ŃL߈П`���Hz ��[T�dZ(R������˛b�>ZC]%&�]�L��ej˃���F�&�-�'��ƴ�y�6yUr;��^-���$;��˚��&�l��jFm�f&��T��CS�:�_����?��w���|�����q�B����^�9q�c�w��ٹ0Ɠ&RAž�'������r^5�/6�#7F���;�_%�R�[Ab���2�drt	�jIuD�9���EF�cb��'�t�ą|�o���fPb���d����X��2 d�Zk�N��Y���7;X��xa<��R����MN7�)ޤ�e�!�NbF^5�Xń����Q�HJDT�����h"�H�`k��?�-�=lȢP�̴w�ۨ�� ���_�>���	Li�UԢ�q���D�[\}~�]Jx
�v�?��}�i��_]@0��I��>_��)JCw���V$��-gOC�P&`*92T��Y�+�º9�'�N�YL٘��Lj�J��_����^_C⁊��`�UH3�o��༄�~y��[�Af��_�� a	g2p̸��Ej,����k�:�vuxF�pK�	�\j�Ω&�[����LW�X4��3�,}x	�ILBkqb���=0$ܒ�.����=Dn���!������}��W%��~(x%��<�n��M��諧3�n��=�G��͔�I\'��j	C�v�ܠ�G�7�`�t������0%¨���#&F݃Rޙ\s�E�
��̾�׽��]Ý�-;C�/��s�����m|�+ʣ�q��w�b!7G���W.��5ꖒ0���k�����֢��љ��i
��E�;�ix�:V�I����ŭ�_�n0O�0�&���A�G拲��3;�qHfN`����P`Y�B�JJr�c6�>,B]�e��EÕlCO��(�p]�!=�SD�� �'�aw�:h &j�R��1�S��c�F�xT��p�,�d/�Q��^��*�5S�a)Q�p�J�LкP.�s	��ZK�N�&$*�Z�oN5/J��KG�a�=�\��Z�!Y5��o=�NB.�\׀�;�x��3����W��<����q2���Ʌ�D����b��X<]�Nyf�T(��u0��Oc��<�A�	Y]�}�+D��sH�R����:�Q!s�!-��Ɔ7q+鐊�*z�t�<t�}��_�@�Trz٭DK��-[^\��"�ya���"�cV[?�ӱWe�N*�����.wJCo:d�h����&OꝪ��:��L�� .���5�K#՚g+l�C_`�a�j�!��de��̘D������;ϴ��;>�ф8c21�;�/�6��s�������K=�$9傎��R4C�;��FΊx���%^��3�;.I
*D�D�_Ŋa�7U�� ��L�<f����V��=�L�k> �@�� ���ۜ������`V߻6��a��:ޗ9Ө���L��	���0i��&�����c�6jB���!��'j��{�R~u�n��8=G�\r5��X|c�s�V�(�%blY���3z�1YH�L��Ez���#Km8�!���qt�!C�&��dhy��8;Y��:�]2��q,Iwֿ��%Q�rr�\>�l�*�)n!$��e��V,�i���ۍ�vC�ѨV�)הgN�j�����q���oHV`�y�T��4b�,ҝ��U�L��*����iKn)�|#-?w���l�o #�!2.�����Ɩ�>]�.ġc%�F !����+�������:r� u"�b�V�M�������A�,b�}P2��� f�P�����m�����T+hx��y[v�{��\ʖqus��d�prƀu��:�/��������T� ���� ·U�r������,� a�^����T� ��|C,��8~S����ƺж�}Ƞ���vۅ�Wyե�O�/c�2���$�82�n��4g�ďMɇܿ���f��Y~}��B��~��������e���ي�|��'�S淙�@O�s��r�[i~X����j�ݷY���gF.���s0��Oŏ�G>�C�.#�S3=��fI��aBn��<�y&�Ѭ����pyY\K4Ȳ0[7l�!�_��Oa	�F9\FޔR�QΔ�?v�h��\1@�P�f|��Y���XL5mx������Y�3�^�ȋ�̴��)�4y5��k���}���J�O��tSe��ר��K����|�Ջ�bPJ� T�
U��}�)��'	҈G���j?t��5o�3�0,&J�,��§�3�N����ҁe�gȘ�ES,�\x*�^�.Ծ$ 9�|�M��|�664@�>�+�O�H�UH6�M�����H$Y6���0�ޫ��;�m��Iho҂��Nd$vAl��8���١�d�K��Yj��^�3ֽ�JO,�8)5��Ek01�A�$��������a����;�bi޽��";1�j�`&����_Vk�p㖱�����yS�������Y�� ���Cϖ23���q&PZ|K��iݡQ�s{�&$9�P��D�I&�!ܛ86T4��<d����[�q���
�LB�T��^$�˵� ͞c���H�Rζ�ϐX�5N@��Wl�HqU�m��.�U*���O��E�Fa����XtBVn�%^���$1�3d24Կc�
�~p�}-Nam'ê�����m�sRy$1�@5(��la�#yd�ߊ�������?m	'�cU7�	�M��a���!�g�̐��Y#�u_�av�U��x�[6��
�ޅm!�'@���vO/��9&/�'z�\K��Q��I8Օ\��Fh��W�`�lv��4��,�����eL�w�.��ߩ[�IC��\�q����O'�v	��:<��K1�]e1y��ICV!���`�.,%����P���p�5�)<�S9`M
,sÍ�y�
Ym7�ͥ:2�����"e.p*L�
fJo�	���}���2���nr(�o��[�fT�h�	l��a�]������K=>�y,�Ŏ�<�
kH4������+��3V��%��rg�%驊��ݠO<;-" ��Qٴ�D�^��C �~�,'���mM\7u2�6�t�	�}�6I6m�I%�7�ZAÚ��\�arr�(�w�֭r����X���@�U�<\6w3����Af�A��BιD�2�x��D�n-��Wbb�SC3���a�������5\�Z}��E��B�T���Gr�ط����S�4:��F�8��nq^�L ����ع��������Y�!���_6�TZB�mMYь	7x#y%�F�w�l��H���7�J�� ���������tҊ���_L��r�92����%��	O8�Zy���N�H�q�	��#?g�J^�#��z>)]�=:X�4���Șd/��
c���^��1�η�����̸~љbje�T�}��T�+ 4o�.�=@@�c���� ���Bb�@"Հ�½����Od��c�`��CC~{@�w*T��g�O�{�����d>��	� �.�6\zi���ȃ0��ȤMmI�����A7G�$�k/jiѓn���Ó��[�oR7���2�W��X� �[`�D�xu�`�7���n��EBǝ�_ �l�9D�~ų���XJ�b���ֵd�Ԕa���u�1`şroK���pk»�Mׄ�tӉ�!����$�/V��9Y���S԰�w1w.0�I��c]/<YD#�����ҙ@p��˦�yO�\�If�T����HM���
9�T%��]�K��.��G(3�iC�v��̞N�H��r�M`�Y��0%���A�Ա��N4s&i4�|���?
�L��e�Aj��Z��.�'Rޡ�C����T�~}�;I1�>!NH.y�i����D/}��b_��������ԷiG�:�Ӌ"M�z<Ge�%u��O����fo���9Vr徆]��=%�tq(3�bb�T��^bc��`�dZ��[��7����>�u�4�B���b�\6�9�8_JB/��t7$�Z�Ow���8���骩Ž�-��<�%z���nPR���3��IjD,�y��U�R�x�2W���
(�=���^S?_R�鳮�{u�]:�MFDە�#����ɗЕ���"o����4/����5!�]�@Bb�sT�)���Pph��}/��,5�ed@)]K������ާ�}l�jb ;�+.N�l��t���&�^qg�~ia߽��5�Z�#G"gj�~�Y���$Fd	b��-� M�j�G�'%���k�X�1���G3z���&�z�ܣ�$t��i>�Oy�h���ѯ�'s��BU'��Ջ* �>��w{���Y��ҩL�T�I��w�
I�F8z��� �LTvL�SL)Β�PY�������,N�#3��z��~I�e��1�0g&W9Mm�	~��?ܲ#++��@��l��@�-	D�&#17��ԃԘ�|��_]S��@�h�I���B���*h@å�!x#C��P���d���ؓ+�[Mw�,��J]qg_z��e�>��)��X�Q��Ea�A[�J������>�^8�|$���#��	'���U�Z���>�ĩ�G��9-KX}V�VV�D�<�{*XMЖX~� 
}:2�P�2�9�9��HM��p�R�z����H������`m��|EB���`��c�i��W?X༘f)(zDC��G���$���>@�;���JVy�	0f�HEe����ީ��)��G�b=R��G��!��*r�v�XG�r�5o�����ix�['�Q� ��B����!�D��H!.4lQN��z-B?g_#���QgY)�"�=Q�3Bk�en��s���{��G��
fF+����U����6��>������UjKD��%W����A6t��&2DA��S�ӯhK�q�Pa��W��]�j��ve��P�<d�-��^ N*M뭜%��1U�>Gێy�$"6"^����@�28F7��_XR*��s5����l��v}v�׋Y�������Y��@��'ZS��u��j@��ҩ����֤sj.ά�X|���f���o����	���ߟ�5�t�)#��oE3�R���LvD=�����ό�'Ɨ%�>i�e���bt��@I*��h�#_� j�Hoѝ�q	P���A���^J �F*4�P��5�"�~$F�!Ғa�$�K���{��c�*�t��z��#�����Pz�-��s��b���J�Pwn�{�����.�� n/�m}�}C 4�N�.��� Cz���p��!�E��=���@�c(er��+yJ��*��V�e.{��_�z�P3�ֹ�M�	`��қ2�*2�G�-(\������_(�.����=���sq��a�	���fC#�d�:��O�D�����p��O�Lވ̜���w;F�/$��Z� I+H^:���������Ҥ,N�NH��Obt[��ѕɀ�HL��%ܹ���\���K���ri��<�ZX��ç*~W��E*�[�{��@�3�4Y�@�J���*jR�Q%v��qՐs{t]��r0W����2@����b@���qd������;r�!�z�W�m4RrG�'SK$.����W0��}x��Ev����w����ŌoE��^F5��g��Tkܞ;L�� ����7 �w{��s�31�h��&=O(�H(~�Y��x�9���F�<v`S,[V�1p�K2#b(��-V��D�[�}BW��iZ���D�f�pe�g�,�~�<L�W�Bx&�Y����L��!G����`\�e��Ȫ&#S��%���r���rC<3�_'9C���'npYޮ�A��X7��3N�m�q���a:9>be��L��RP�ww�_�d)Is�p*�i�j��я�Yj%�D���is
�A�nY����L8��"��Jj��ƶ�%[~۬Q�t�����K��C���������ol|�_�'~��A[~�d�t��C9�_�xY#M���' r���g�/�|
R��<މ=}�Q��j�L|C�A��u��i�c�L-Y�������wfy?a�o#� I�N�%6$'7�� �]�ͣ_��gmz���9�ݳ�6�wW|m�g�NL��|��yP�ۆ���-�|Zr��q���C)
��Ԍ̄�jC��݁�n)PU�6'@�3:f��$Խ�k��oI�&93�|�p�ĉ5�񠦍\JP����+|��h\�0�$�kҶ�jP)�w�ze��n���Ғo�Av���ѐgh��k��}�{[EZ���{�N�V��y�G���X�Э��	iN����d�[HX�yfCPl��qQ�@@ ��J	��wp:����� ��%��ЀoL�3�$������$�d�I_�~Ǳ�y$���E��{^SL����~���YihN�ۃO�V��r��6�"�Y���yP�aR��)ֿ��޿��(�Xw�ZN�d�o�jx8Um��[�e+c�o�"yݟB���x�Y39ȏ
����-i�]�'����NQވA�fЃܽBx#�g���(p�	����63uv��:*��h��7������낷����J��4�
ݢ�!��[�bv�54��Ī�{+1�l@];@���v9[�
������Yk�Q��P.�%H� ��-@��b����v���i?.Y	!q���A�,��`�Z9
P3���}����r�k�yP�'��%�$:V+G�Ȑ�3��X����ӯ�d����n��/�0���FSZ�=�V�m���nI�_���2��%z��7Xϡ����l�/�0`yd�eI&s�!3�Z�N���q��l�L<�/��T��ٌJixp#����U�i�[����v��:�=%�c�-#Q֥a�h�*�Xy��}6�{��6.V_w��D������r=~^��vz��~q�Ⲇ�#n�#�w�%Z�!r�v��g^�V�����I|��NG�d@"�%1Ag|�C�]��^]�$�mu�g��E@�GRiJn�����#�z��@�_ϴ\�e�mσ����Xd���
j��y�2=�:5���o�����M�'� ����G���xJ,���g����*ndR��bE��a:������&�0��Y���n,�J��ŗ@����:o4,1�Mp)b@�خꆙ�$}u@���m�-��}�-u���=��G�����7x#�}�xt���4�8Ak$	��ꪒ�<���i��Rr�]�Ud���7ā�ؼ_0AR��*Lܐ�Zi�6ו�쨀�Q�_����:��︇��o���q���0�t�x��pS�(�by7�ã�)�8Q���l��H��dѽ��� ӫ'��I��򌄰��F�Ӟj��g��F���Ȥ_��G>`�J�㜁"��4����# kUL���:�O����Gn󔠏O{]Ee}�����6�M��iV{�c�%�1����CZ�(^��`���)T�}j�6��q�)���!d�KU��c����V�yj&9R���x���[7��n�f�0?�
�Q��og��y��̙�D�G�J0����Q��aO��K��N�yf�!	^��Fb�ַ���ѻ��^I����d�y�Y��t` !��������+���D*�_c��p��
VDFJ�*�pGI�Q#�4�[���u����ٕXF*�x�:a}e�`n���_�t J�NH���ڟ1��TΡ���s�m�DV��9be���q�H<����k���eݱ0����u�T�y1�����w�[s(<>|B
�rQ��ٴx��l�O=9��X��oT-˕�%�lz�-��@C��1��g����3��z�E��;UZ$��Z�ߧp}E��. ��I�:��9����E��b��};'2m�z�lQY-D�]���A�/#��$4���xg�}0�]�.����V#��M��u@��?t����g�&�{"Ր���]�1�������L��0�s�W}p���k_�'��`��yN99=.kW��d˙���[��N�E�=61y���s�f�Ր�'{%ҁB��x�B���S��w#�}��q�>u��w���uAG��s�3�uX���:����VE������ಟ����`��W��_,����YK��Fϙ�e��?���ct�����]]����d����樬��k*T�&vܟ�!�=�8�S\|���˳�o�'�5Jm�sj���~��9�hN_y�t��w֯��?Y�j��B��HS��KZ���D� -z��4w�P,��*�M\���B�@l���1�e������ު���53�*��#;����R�:�4��rI{�ѯp����3�3�}�b�&�λQva*(�Sq,k���*�gh�գ�ۏ���_Nu��8����������y��V�� '��Uy�/�G�V|6%@�1{�w�k��R/u*e��)��Z��W}�r�kcHx�M�bN�h�L���W�\ు�ޜ���C�.5Ga+Q3�Vɏ�(�ǽpǡs����+8¿tf�"w�����̟9RJ�O��G�~��m�|Z��	tS��`�����z��Q2u��yC�Pd���<o�~^�V�e!�4+�Ɖ�OE~Z��eJ�p�!�K��~��fv(�R�#(��e�����d�~�lր�Ė��׭�H��nHVo�P'Ot㛁��\�f���b����{�搴�š��p+Os�&�%j�T��Ҕ'Ɩ���1�'(����/Q�@�J(����]S��w6o�v�{�I �����^�K'��k��ǂ��E�D������F
���?�̿��L�P�e��.2���zn&���Ը�$��v�t\F��MF���	z�]�{N��co&�B&����P'�� ���i$4�j(�1-S��j{9���3T��%l��f2&Z����͝�ԙ��YM�*^��������.k�s�9wr.}�ZS��9<�k<��z�M~˯ �p�f)�ݴw���P'*��=��F����0��j�頉T�r�Y;�Gm�D֕�b���5�ۑ���V[�A��E��{3���2�I���h6�o���=ᠷ	'�@��twZ>�7�r�k�gg�z͑�'�Nr%�0���=�+������є��OM�n~�R�[�
zFH���C#b�e;e�vYyT�d�2qk�m�|�!�22��5n��Æ%5��h�\Zצ��z��fW*�*���G�M�X�M���9X��w)�6V��S)���aݩp_����)Rg�Ǖ���	^��m���&�B�í��^�:�T�W|vAU���j�w$Zo7ᴥ�;/U��i����uG����2���`O��vQKIr�y�A �ͩ����ܝԀd,�6.�����ȓ ��|�7�"�H�P��ѝ�)���9Ԫ�������|~��b�x'X�M�igQ��^F��I	�{ m���ϗ?[k�V@��.X��قE��O�#��_aN7��M4L���fj�0�M-�hp싟��s������(��=7��޳�j�%NGT�[�����J�{�7	����4���:�1��z1�_�.�˓F��;�7J����
�;z�����*�k��t���lM�V��Y�+cآ��%��������ӈ� !Ҧ�p��_�`*�� �>����q�>�k�<cˑ �o� ye�������HfNT��(��ՙ�6E<�"�<�f�p6�:��.��5�����'I��b����5,A#!U�����P���inu������?|��L���{��.=��] H��Ju������W:|� ˪�z��5�n�V�.\�P阎ɸ�%������l4#G-��n�מ)j�r"P�tӚ[��k�uW]��d�T7�3��.Cu��7Nj}�.�e鲪�&�CF�b���Ќ���̏��^��f�Bo=����	j%���e<z�gf67�F���A��ԇ+e}� Ф8��m��ٓ�3���+������ZQ�c��T-�&X���_��*ϊT��J<YA�u
���N�ΔԾ43z�+T#U��d�~���(�RVY��}����^u�If��\_��Z'�LVB�� ��,�|γ������Ø�a��bV�P���X!���hWO�A㦝w�����b
oH�h�h��p&�[ ��Mb@�g�UhiZ\���$r�q�^F��b?y�$o�1iQh�"�.���q�}��
�����Y�Q��:Ze�,�;h^2��(�?�����iτ<M&��^�A"�ɏ�G�jnM�߫hR(+|i�����yN_Zٔ2�6�5�j���x�DO���k��>�g��V��#s��'�h��Oy*خd>Y� ���wѫE6�aF�w����/���M=�KGÍ�k3�ϓ5���N_�P
[��e���6��K��7a0#d#`g�G>��O�9H���_�)��MCw���bئJ�mCZ�T�^�^�<x7"c)3B�-i~����I":v��T*أT!�m�o�$���� ��x��R>Dː-Bg	�?� ~2�zQ=Y�K�v��A���$΍���z�%��B��ѐX�E�.���*��֑�
ȗ�M��rPUH��ȅo��Y�~`P���t+C<q�� G�7,A��I��w �\bWg���6��K8�*��C?n*�)�Yix��0�S��L�����[,$=/#_��/(���L�38r����V���y*��М;~�m��P|KjgjSCE�Ȫ�]\s&=h�81j����:{`���`,q%Υ��P���hP���uv*1ۧͼÔ(��C�;����5�sN����F�Cғ�+6�4����Cƻ������ �mئH���W{})�iO�>�ݰ�RI�t90ԫQ�3L�?�)���}X;�8ð��z�g3� �����z�I����עb\�R�>�@�c��(���A	P-��sp��QS^��� 0:|X�óL���V��S^1���G��Y���7U\�̮�ׂ����Vo�W�cI�ǍY�kU?c��R��0���r��/��؂��$�HuQ>�3�����g�;�	4+�J���
8/�|'e��5%.�o;oa���{fa"� �oLn�W��̍�����F5�]!HP�!�+wb��:A	d�%f�(�iG{L)�![��>��"al�P������<_ˍ^����c�/I�fhb_��v�k�����B_i�Ƭ�|"��g�?3�`N�ex�<����dq��BH��f���G�c�����J��
��%�KZ���^H�}�c�X�^:��˔�&o���zڔu����c��y5���LM��r�B��P����qt�Б%�A��[�������P��,�G�9�R��ff+�� �U9mJ,��y�f��D�y���򮳼�
k�K�a�'z�~]��;�����U�������@	�������ʉ�P�.�ƹ���#%��矦�c�ɵ9�\Ȣ��F��%�~F���zU
���#��6M��hq��oR����W�֭��1� �8x��r8&S�3�Ml��-�|��y�i�Ʋm"��<@窡�Ax�#+��6���_�h����T�8���������9�r��"J�����aOt�p���9��e���g>����4t�B	��j�`CI�(+:=��=�w�/����1S��p�z,Ma%�ȝ!�}����/���E(<&T}k�z�z-'˩�zO; �ȥ��(z*"��.=O��Ӎ'��Kށ0�������4�Y����i�����?=��-Ha�� �+4& �h��01p��˲̣yk#7,��^��@/�����0e��[LBm���ÔM�`��@��!nW��{}�_=pn��v%�T�B�������	�gz$����vu�+���.�;�"�ʎY�QBc����=��6�MG�*@�o�������g�cɲ^(��d���R\�Dz���g��a�cU}j"��{��4�i>�V,3�V��V�`>.@�(A$�C�"]Q�]O̥^�w|�YRW��"Y�D�\�W��sH:���)w�����`+��4��8����.T��/'<��Aol���|����Lr��d�P�ٍ46���Qh�l:%�R�l�����5�nI��VwSP�.��l�m�KVc5D�b%a_�j��Fi�@1�_z�"��S��L\sa\����4��bP������y���������Z�:��#�i�T�+Tڈ;XX��i����V�02]ͱ���rg-�=w�gH/ ��"dѺ|h�d�p������9X&��<)��9�+?{[ �M��1���Bt>�1�J�$�'DrÊ���0�&�?�_I�%�o03���k"����s|ټ�����1�(�\B�]]��Y�7F�fR+}��݇�y<�I	_5����`!�@��2eE<X���G�r2�}x�Xu�X����T[�nQz���Y/�-,eo���n�Z�kU���d
��:��X�[�8g�SG�=�Р���Mi�@��=�ꨰ��<�����Y�l�/�mϷ���D�k��^zo��E�L�V�
͖ND~�	=n-;"�O���GM"�t���c�<��6}���m�s�Ѡ�[�>�4��غ��s��p4^�H��[�Խ�X�g�G ����/��)��;+p�^�%J[:q�����^&#}.�U(]�Ά.�+F�����ܫ��1�]G�/�D��B�c�p��m#����Z1k0�|��Oɽ�(;g�RP�X��/^R���X�����%������̀��5�y���d0�:\w�AVI*A��5�����#�		����_6
����8x��oE�	�IH����}=���jn��k֠̐Ql�鬚�+E���uhr�P$�-00$X���W܁�L�wѬDs�oq��5��`���)� |zTχb/b4K�:m�r{�¯���Dnh9Rk����3�z|�S�����Wo���)bEvH0��7�H4�k��]�?~Q�%�d�T�}�@Jw[�B�����޸���䦙�\�Y�͌�4G#(@������y����hn�.�����[@!�Չ_��
(hZ� Y7�-R�U��?�Tv���+���`����_:�����vT~���3��|J�zmM si5]�1)�C�,�,��,@��!�N7������	眶��b/��Q����1��9�u������y�cj�>k�Lh�R
;����ګ��[��Cޱd�,$��ry����)��eg*��/͟W��M�.�#`n�J�EuO��~�f�|�#� ]�g��?� ��>�e��7�4��֟�A�T�9/U裃}�j�
��~橆��P=r����R�O�Z(��?uM-�* 1N��x��" �q�6��&���]\��>�$η���.�4��C+ݝ$J��Hl!�m銛g�j"K���W�Q�1��K"�\��3�om/P:����t��΀u�v� 0�����"�Rd�������wKC��lg�Fƀ
��lհ�����x�$��L����W�S�ͤ�|�u���)J�B�dh���kT� ▐���Ȫ��U)Xd��ňW0�94��=�3�y��_�?'�	�?ku}�q���ȋ�!�ڼ4�l�ye}�qC<�}�ݶ�P[!.n�Ybm1(T	��jh@}��=DU�
�7A]���J\x�h鹿�)����.NRqX��k���n]���l��Zˣ���SC7�< e2��s�ڔ�⌂��������4��6�$�8k�K�޻	�.e��e�Eް��!ɍ�#2������x6�ʿ�����ٜy��dT5�p��~��6�)- ��  1F%<���τkN���Mv����9`%#��S 8a!ӂ��6�9��Ut�I��`w=���\:'٣�L4��Sf�{%oo�-�6ㆨ��A2,�x'��ZL�����O��k�´��$������@�ק�j�����H�9�ӾY)��/�c yĽ�"�7@��ajE�'i5������{\e�k+=?kF���3O�U�,��
&���;EΓ����a�uj8l��C�Y�GO OaU���z��x��F*��D���icj8s&��# J@C���
#�N���_d��)`u���zΟ* ��,�B�!;��t��"ct@4rrZd������G�5�P�O�ۿ��z:Ϧ�Vz+����=���fK8����֘�
���8�,��s��9��HuRB�Y�C��p������&iC�XD����X�d��P�Y�X�;���H�;�G�^�֣�P�����Bi'��%�F�L[�u
⮁�ib��<�%`^����'���=1bx�h��
�a�3�I�����ӻ��저�	,��mHzb�{�*H�Vx���&;(��-�	KT�x��۶�p�ϛ�2�RZ|�?��y��ES��q�P~K�H�$��\�����r��dL�E=S��ق��ɜo]�訓�!,�X��x!P$�1!E;5ɵTs��pZU��R*�^�00hϞ� ػ �,y�B���r|[]��<[�{�͂H�u�[�&i�X������	�Z�
Kẍ3�k�1����Rs
����]���v,���:�?{S���ω�����H��|��%�x(6�z�9x�p�W���y6.%�2Y�f���]�c��)���>�dď ���:ye�r$�EAЦn�Tq窆���|���I�K�(m��5�����E3���@�0��}��@�J��2��rؼ�ђ�ѻ��Mt��e<	 )��Z~��F���?�&u'gK>eq�:`O�T��q������4>NX�u��/�X� �\^t��GM���h�Z�
?������~��C5���f2n�c��~�X| ��N�Q0��F4o�!H���YG06j1��Hq������??D?g�(h�b�2j58([�̿a���U����<H����Nq7��;+n� ��A��������,�P�2���k䒴��}��F1N�{�A�M��4�=�܋�ŷ训([*G[d�H�`�}ÜF���<P�YH��`�G����?����Qx�/8֞E5�ev��	�Q�_��|�D!�7c����B���3��i����֒ �0����#zR���6�L?gó��Ѥ�ޠ�����L�Q���=m��<�Z���=餔쁌��P@��SrAҹ7L=�5�W��9k�&�&�$�+q|Y3�ť�DJF���IJ:K�LJ�P}Md�C��e�<Я-Wn�ٔ��3�I��P�T�eb�/*s��BLn����-�+GyNp�M���$�_DGb>ݱ�k���Ͱe��ߟVo�GqLe��i�P�+@�	�##�r��	�(Օ�Y���͌v�Ku��v��MF[ �z��j�_q9AB91(�"�1F��[c�7�F���\�?[��o�n�d:��o��䪚������؎g�&��Y27���8�{�mW�k���_E�r����g	�2����A�e
�,$���MI�|^��������o�[NK���'��Jp�.Sz �L�?�߀����02��x9�Fl�-�]S���O����Mnk�sj�SAº��(�JB꬇ا��څƗm�2���8�B�57n������Ą�L%�cg!��D)�Y��|��7v�8��ֱX��4f���ͤב���P��mn��\OJ�I��w�^:��"H��}�k�����4E�ӿem�%4��j�A��L�&?ߎ�49����}��$�sc �S�'-��/9O>�X.�::hBK��.�Ia����j�:$�a&�?DVI<+�J�v<`�U���:�c0��
s��ç% �9�b�ۆ
P!*����s�~�p�33��0 g���`Y�z;��$�|��A��lh>Ѹܤ7��r8�C��G�q�D�跔�� G�޸�gEw��^E(�4�E����#�?�~d���|׷��a��H�!'��$����h��g���.`�v]PQ�r�hﺽ�m���f���#b����蔃�!s�l��O������n��4͏y�K���m�����sYyFh������PU|A�i�YX�G�SÚ��$��8�̈�IR�-eON�mf����.���I0�
^{���3�%͑&+S�,��%0�s�0�+E{a�A���/���0Z)������$�9�|�Z?��Mk������\��>-���	���.Mk���R$�+g�k﷾a&�
�Ɯ:T4g�ꯊ�3?�2]7u�iC1��+�|�����N,�YH�y,�
Kɭ_m�E����!�	p��=�TMO��ì�p�f�5H�^*S\��D͘�M�c���ߔ7��Wfi���Q�������n� %^���Q�'�p��2�>Ґw���vf �����\*�r��x�m��r�@�M���o{\i���p��|�M-X�'�K���"~���
ά�W4~�$z�	�gƙ'a�G��E;�̨�C��:�s����Sb�n�ZVH ɖ��g��v�*��m���(�^ʝ`�
��~e�Asa@N�W��h�&@��KO&y9�a˺�M��,1��%��
P��:�FP��ZG�Ų���C�h��H$���H��	BqI�ۨ_���%Z�S�����2Eə����ư��/�I0�?]$��%�g_7F�c��E�f>��/ݺ��Ϩ6��?��=7+^E��~��B�)��X����
'T'"O�aƧ���A�fS�^�Y�+����;'�@{f�"��Q��P8Hp��s�M �[e�`�_6r�����ty�~1+؄�P�zU�$���WG�����[���'��a�eШ_��ln���+�B����q�ۮSo�f!���ڣ����f�ϴP�r�������:�H�r垯B Ȏ��$ '�{��]ta-�����b�5���Ls��6v���홬_�$;�<��b����f�khD�mo��V� �4T�{ą��R�ˉ��~'"�ԯQ�U��N�
z�#�ʅn�Ӥ���o�>�gX9�91㫬kb�^�eb�u���D=�Gg
0h� ���#c�(�D=k1?�R��+t7�I�p����P!lIW+ݛ�#L����"x��#D�G�psj�1)�Ygj"�'�Û�F��O�Z�oqLC7����n�㙩EF�O�c8��p��|�W��B�����@��ءp08$|���Κ\L����� ��	�Ql�Dq.�0�h(���j�+wXt�/t�Wx�Ii�즏U
�/�� ��:������qK]Jm���Z}$�n�
1��%�Ԡ�F� ~s6�ˊo�<N���M2�v��C�nEdm	$�=�F�]R�:+-�=0�V�"H0��;`v�7��8�҇�� ��i_[����c~�7֐ǳ �ET�V�6��9�Eh�
�KA�e���nM��^$�n��\�$C�$��ɐ�.���+�޴P�&Oś�8�~��ȴ\ڕ��~�%�qn�F�k�O��|�m�=�`?Et��
�Z�H��}H�^�ck�sg\'����4�B���h._�x"�d�NL�$طؓu�D-�RDN�#�m��k(��4�Q����btW1�K�@L�X�7�����;�E���
ѩ�����~��x�f�j�`�F��Ή���)�_ ؒL�Se`+G}`A��x&��c��T�%29����}��&������ậ�F^|ޚo��K$r�w�A�tρ�O��А�WE�#&�g��8�%Éx���(GP��Y7�ǌM2�aaK2=�nh<y��+�2mZm�7.?8<�\V�Uvش���o�L���=���d)Y����&��Wñ��|ˌ�΁BX�/&��yY��� 8���`K�x�V���N��������~߶K��@yz�w�"�r���%_�����p��V�u�{l��o�)�-��z0���=��a�QzqV�Z���z+vܜ�X�&PH��%���!c�+}���S�Y�`��!'�|�J�=�jҴx��\�2�c o��|�9�}j�;&󄁲Y�}#��ke]A#�[H�]�g,�n=)��A	e�P>
:�ԇ�J��z�h�"����n�M�ܓDn&��hX�_���v�%�&7�>�kj����K�u�2�����c�g��ۇ���
Q�e8\�ػ��R�z�����scor�&��wd��Yp���0�� x�M�*G/��6`� 9Z�U_�t�����}�i�A���"��tm�Bٸ=��t�(���u�eՂj�x���zS���0����nx�v��N�Kb��J��n���#S���X�����o-@�=I�(�*&�fi��ʐſT�r~|M�f�&z�3R}������2O ���;��QC9H�j߂R֔���s���SX��A0̻u���'�;�2Reˮ)I�������P��uc1��oЂ%z�l�=��Z�攤�fk�̧b��?�2�p�[��J���t���^���Jݗ+̿����h `��d�����h���%�g~����X�w:�_@�oB��^w\fPO_�S
aJ��+�X�:ٳ�8v����Ɩ4d��&�t^��{���l�b��7�R{~9�����Q&F���vP�'�Ϻz^+�a,D�����+<#�����u�&�c�;	6r�j)��Ɣh�O/bۤЄ����d[]2�N�$B���A�b�ޘ����#���ߚ����������	A�Z�u�6GJ�46�W������ј7�b�������w :j@���o��O���;��έp ���B�8
A+8��u�ɭ�#F����i��G��
���Y��Z���>�LVF7ڭ.��P����3Fd���H�9F�4��Q��)�\6b���\�eG�V=�!��?B����e�R\�dT�d����-�e����J'��7�_�������Q���iѵi�pUr_����@�½�.�.%7m
��\A�"O��bP��;YmW2�r�fz�HB��0=���L]s2����v.4d�9Q�j�`[���S���(@��XV
�.�v��zJ˞/�����ă�+a_g�a����U�!��
��%(���Ieh6z�4+�(u�29��vgvc����4��.(��c>�l0����ڵT�0�|,4U�|�w'>"��P#ġ�xB)oA�%H�Dm9�M�aM �U�d��4�{fY����bU��玊=��J�Ct�|�*U�Ǆ*�в�����R��'i�2?���I��&s�Ͽk�}4�j�Z�@�V�%x�́����cJT�o����8���Z=7kC�a���*���=&]��b���pS�zE����nݜ��?������m�B'r�_�rx�P�2^h�o����,��˫?���+OG��4���Z:���kg�BOc��y���F)��]
|MK2A��z9>��-�.�?܂һߺA�z���AI0�uQ(���M.l����\�/n�9�D�%~g�r܉~Y�������5	!�B���8h�P��ms�S[63�h�B{,��%E=p�'��b��`\Be�I���?�41Ľ����Z�n����A{2��HF�HLϘچ{ې��k��5\�ɋ�nQhF�Uf��ч��.�6PG{�plP9��h1|�H\�+c�$Dc�����m�y[��l��Mfv`ʯEa#N:�W ����~a�4�����0�P��k\.mqV����r�u%뿭� 6M�#_�b�R��m�ڢ0�+�ͅ�`�o����3OBk�������b�����l����3���nQ�{e6��Q�J\毅
�<�L����ho�9�G�A�s���9�2���Ai¤ ��h�{N By�Z�B(�
��v_��1�(g[*�>|�<9��k�W��3f��Q/!G����1��CQ�
A	�G�)=*SQ���N~���|�Yv�t]5����~T�V�咑��~��ٚThaz�(�5IR�\?�g��}W��^�m�:�%~8P���{���a��b{ &���T`���Q"&c�ة��,�93F�;^�c�E�������A�b<�47\
��z�j�������&���?�4�?������^U�Q��3��L�w�Vs��V�g�,�,7*�E���PW�������ܓ��� v�ٟ1mzJK�BNeBǁ�H���Ĕ{�r��� ��5�����ν��q_��-��m��/$l�m5T��C�� :`X�58� "��)X
�����\J��Ԣ{�қa�}/��Y�I�8(	�D"�rkվ ;������N�a��Ц&z��(���<� o��E��@��$��_�0kgk�A��r�!5��?��34����zr~,��W��m�$����� �򞧉�9ļ�b��Q�r]��Z�4%��Y���?-lv�6��߳$P�
����ٽ�M�y���bt�73{�=j��q�~����MRɄS����+��7�B��( ̭��'1�Cj����Y�S\�x�r��~�"#�Ctt1a��?7�K�z�u3��I7�-
��JܜcDM}&(X�A5>������3.�E��͂Şf�p��l�����Y��)G,P�}�o����+�y5HQ����!����l� ��@�*��I�|�'^b�d@���R��A�D�E���aX���cO�'�E��_�ؼ$��`��ܽ�C2%|�JXj=��::��R<��+�4�Վ`ȉ����I/]x`�9] n&Ƣ�ڠ BT�MߪuU���9 6��I�_,����f-�����bd�C���`��ep����ʀ#�e'�S����!=���(r�װ��g5����������O����NA����T�y��¦�^�ݡ�ا!W�pE���U�|G��`R3*✙����h�	&��we)�6��/ږ�Rp�V)(~�$пY����h�!N�[(��z?���[b��;<O録���Q��I�}07�ZWϓ����Cw�w�av�S��=�%4�QR�0aK~�t8�H�.J�{�Ʋ�^�
���Lg��Q�+���0I�2��ۦ�1	�Ah�ƱD�b��|�?E�V�k�4�{�ci�5�����(��T��G�S�C�v�}���ͪ��#�u��/_�[�#{���3�ѯj�̲	���(�h2%�}8Ȃ{��cu��d�`!�d��n�-���-��+���.=R��F��-n��?�����	�7eCs$lzV���\9P���D�p�F�`����.�S}eky�]+uI:6�M4�6U2���K��O� 0p��X�]ms.QI9k������O�����i�t���r�^��_z��IJ��=?�=�@��φ lͶ����BI[�6dR�����z�נސ��,�~s&���q�TZ:Q�]�.V�\r�� �n�N.�y���?mG0d;��Zm(�yF������� ��:	l3��-}Ha\Q��5��6 �<.V�LlԕVT���}�Z���<\k�@����\C[!���T`�r����:�Vn �U���q^�B<a��Y=�o8l ��h3�<���i�D�� ט�����{���^�E��KJ�&o��g,��yt'����Hf�qD���b�\��9��+]?�U��`�t�~��$���z��=#N�C)J/���qZ� �|��w�4���������A�U�Q�>gh��7�O��"�~�K�Н��
��i�r3n~6	�s�y��0b�Zc��m��d�h�^e^U\4�\Ր���ԅ]mj�]ex������1�[戼��\{W4�|����-�#F�Ъ����5�E�45�-xLk�c�gL����W� .�V/X�(]'+���S��[Wؕ�8���T���-z�!B^jI�*��K�/<��H�ߊ
�ax.0)$B%�+@��j���n��F�k�
?��a�������W���l�5�QP:<��q�����k�H7���d���7�@Ӓ����;M�<�M'��z��f��I�g��ZQW�\,">Qd`�+O?�^4;�2$Y�����q�W>wςh�-���s�#wuu�fn}²G��k�D����7ȰF��⡗ų�����D��X��ں�&�i�;�ķu4���jq���ŹV#E��0ᡣ�6�2��'F���u����ӓ"�G$F$�ق��J��O�`5�%4e��U��ӻE-$B�L�	���J"_��I[ul��&��m��<A�����ɇ�#:GC93����DWP����]N�ɭ]ꅌ(�f�=��8��m��ܳRs�N;Ս�m�И�8�����hҊh����|���t�⸓U�����������QZ���d^�4B�Z�F%����TN��Y����b!7�d6��@hx~���b��}�k�P`u ��D,��n_�B�t$��:g/!�2��	�P���wRΌ�V�o7ʫ�0�S��մ��K�Z�p����L��y�:��3IVѴb����P�hI�\�vu�x#i����\�eI�(�٘%���9��	唫��"b�C	�9f��F��U*a��؂igQ�,A��:)��V��Sb�Uv٣4�6�0I>11t��P'�y,�K���Y7)������+�ؗ�'*Q���oI;������#vQLF]Ę��ͱ+阍3_7�N���8�f �؄�O��'Z����pMCR����<P�D�DW���#m��� �}���e�oT��b���G��E�9߇P~��r�_~#���H�(:�*	*93z{�4���!���۳g���@@}m����3=)|pܗ�W�����[EP�O��⛒t���Y�N� �)^�BwC�UOe����].K^���^��y7�hZ�)@�OT�ޘ�kL�Ѹ�HT�l�U�V����"LP�}/ ʻ��B��7!?����k�JS��@��If��H�?��.���sE�����i~��L�Ě�r�����d�cIi1��nl
��YB�]rG�5^C�ί�}8��%de���	�L�����L٩�n���Vc���Q~�"���evxX����Mays ��7�qf�;(�;��I㐸cD~�m`��u����(ŉ��68a�S#��A+���FDo�3�|ثb�)PSnH��g=��Zt�j��пɣ���!J��$7/]��8$�k7f	��U>6L	��>j��~+b 
�Z�K����A���j�������g��&����z�,����]\L�~��Z��>�n����{l����w���M�����c�B��$K�z��!B�Sh"~����D��(Z6�=Up,aO�}~fˌ,�g���u����,g���e������*ۗ�Ұ�\^���N7d���	}w��rrm�~�)��)�4v��װ��axn ���x�<�����R.t���Z�O�j���?��냐(����	2~�:*� ���m4�,~��!����B�\�!%>�Ucލ��!#>#=hO�Je������yu�.���O��/��Lj�$�N���xmV�&zx(�V[$-�w�X�k��'�JIrCH���P��V�L�߻��޺BH�ξTM��WZmF)m��5f	V���> N퓉v�	[Q����[oN���!w%'��,��0�}��>��WYָi�iff;/��?�j�{���V�Y��#y8��s�c7�Ӂ��ヘ�t5*�s��cxbȀ�x[\�z�Т[�4�+3 �^���D'�W���W��KNL�]��Au���fؾ����6�`	Su?�3}����O�R�"><(��2I�So��Օ
��Fi���?��^��ro�ޖIz)�$ԇ㟩��)����c���8%I4Ŕ�cEC��86Y��ox�/5J��gؾ|(��{��m��Qn�jgo��� �R��mftW(�D#"<��Z��}�΢H�)n2}�*��Pv��DЖp�B�j]�SM�&�8��9�n��n�'�.g�$�	�@�9������1��p{nw�[��Ҥ.F��,q��q�p��]a`O���^l	����Hm⒈�Is����9��Ꞛ��c0ʞ�C�>�ݨ�m��&��
ЕU+äG���bz�[�#F^��&�?��u��68��4�m]Ud�`�5	ԟ�D�-Xr�;o�����X�0��W#8�vR(7�ot�ݽq:7ݟJ�?U2\L��I�򁯴^��ܪ��
���>0ӱBhp�R6+�H��g��AY�BV"�T̺hO��bv�+L��z�M֯I�`&<�C����iY� OOӇ���*��� ��{��x��g_q�AP�^
K��-��p����k/��Q���̟��F���*-�c>���ma�N
�@h�mLI�<�kG6/�
�C��)ܥ	� �#i��+ ��iNco���<T�c]��.��(�sb��}�U�6� ַ���O��5L�6�b��n�?q�Ķ.k�]J`�G��1���ߞ���^j����VZoob/"z4����]��q�ih��׆?6@�10 ���m�J"A'+GIA{�r�0[i zT���!�����"�8_�ZN2�0�W���D���!�1��||Q	+C�ޝ��(T�e����0\}+�3G�}-� �OT�:-z���\�rD<���pJn�A��ߵ-5���V�~G��wB_�E1\z�\�+�BāYܶ�vg5��8<i@,A��s�{���y5�:�f��60�Wx�7��/R��o�Ϸe���\�шw�>}�	��L������N-����?OA��!��Ǚ�?�w�U1b$W�����W\1��]V�z��&+���6J9���w+���:+>U�&y�~<ԒѦ�v2Y�����U�ú��ˑKNm^��|��V�q��7$o���)BG^�ɠ�n�#�ϴ��Pb]ݔL(<�Nnӕ��L��(��J	��8#aߣ"`�v��nYϯq����2��R4�ѕ��0�׌��qVD�1rp�wtzAď}o ���F��Ï� �5T�]"��OV��SM<�F�-�o<����C��8����ݶo�{~EsU�����<�E�8�k����}�{̈0қ|p�K�g��ѰA���sX�.��d:-nx��͌m���D/Q|�Bi6���+��쥒SO$!�� ��Ò�Brk�L��j�P���VW0B�MY�p2B����3}��7<X���F����s�k�b��<���H-�����ج8���}��b&D�q�'R�}�R
�����/R+�J
�dc]�����]� ��Y�RU ���9�D�3=�=��sUT�Z�gιƁ�B�3��^i��2�����`�@�|��k!1yB,ܠ�JF�{X�ۄ����oS�����Oj�"�P� ~w���v����5L?;������8l5?���T�F��b��D��j�6���2[���YǛ	����e;��"*�57� �}�p̐Ә����l�Ʒq�p���&٠_G�!]I�z#>���Hf1��O����f�K?��A�5�j��si	̀�oA�5�D[��ذ+���}�{E�6G����ߩ�A�e�Ţ�Q�r��f_FEi�Q<￀wn�Ľ��g&�j���B�hZ�/
�iA��co[���P�ūQ�� �Y�y6+��b�-��B���N�؀r�ę�d���n��ς��r ��X9�>�#Po��\�k�����m��?�'T'clEa׭�ε�U_�x���=��R����o��*�z�1ɈEG����+�L��B�g0��]�oD�ߪ��qϩg̮�ŗ�wHx�q[����ԉ{�q�p���_��4�.�N޷��WZ:�4Q�Ys7����}4c馏L?�=Y�&ƭ4��aMR��n�`j�ݮ�Bh�sO��6���NX�Ϫ�LN]D{�DE3{�e�&Q�u �=ɕ�+ugXr�\T}�����8�ĵD��r
B��ؐzH� Fx�,����܁�R:~���J�ݿ�Ϙ.��Z!�gv	�oX�Ϣ����� ����}��և�?j4��!MM��#@ �q�g~�QP�鑑^���_�敲���f���q���XMO��UW
�x���.�����#&
�bM��CU 2�Pg{.f����)F��T�P���IÓ����7Ϸ�pzTl�P��n^~�tN�m�Qw�eY[��R�<`��_S��mX� ��rڻ��ux���=�8�"��tB3�c�3[מּ��t0��4	��j�9����RK�P����R�(����mE�׳�w�ZXS8z��|9,U��ѣ�/�p"��4-���Oy�LCGe��ԁ ����"�H���@�g�%W��;�(xt&8��⌭(���"�����G�5=�5/5~�=��8��JU2����r
�F�4M��$ɞ�����Hf��os2��n�3�H��c�KXQT ��]4UIES��j�?�#�;|Q+�U����y_����G�U�</}�ޫe�|p��-TwF}�~�l�'z�*S,9cR9���&��p�ϩ���R���'W&7�ۜ�H,t��*9�<�Gĩy��EDM�2���r�Is�ڏH��^�B�m+��c`��������?mNEU����|�h�t����E���y�q|/(��%ʐG6���3��JQ����y�����`&j	Jhc9'�:	�#�*��.~���7����kƣ4
�����g���1)AA��]Ҩpq���3�
�,�����P=?��	��?Z�MJ��%�]��Y�=8�cq��fo�W�b���~�}z==��/�aה��Ƹ���%PbHc�W�6��߲`���L\��n�a#Zͥz,$��_#h�Dn�@����\��\��b��M��,�+�CJ�~O+����³M�F��Ϧ0�kx�8�mJ4ɺX��ߊ�ڽ��!̚��~�P&K����1��	�<U
�auNGx��Pl�XR�#N3$r`F����Z�'��_?��/3�o�~��&���*�sO?���(/G�]�����ű�ES����\ߘ�G�w�-b�K�?��a|9�M�����;���[���W�\�s>�r�M^9������ٛ!d�BTQ���h��T�vO��yu�#{6`��lzi���P�����Ai OW�����,D*���t�ן-�DG^�ʏ���˸"��7�CXI�0S�kf#�w㩱�/`4	x������ńC�|��蠐��|�1��3w���[Gd�?K�U"���
������lh�O]��?6Z����Y_��X�7H�{h�h�g���F���� �ho�$~�<���ܭ�����q&�n]&J=A��%a�$����63�зTj�vk�,�A4�aC�����D�Hk�Y@v�YW�c`Y?[x1���/�w�2Н�y�j)(�_)�0��������kB��z�t�e�/
�W���`�tB���6�?��O�VS�)�Y����{��L�d���y�x��OY�:��ƨ�g<g'�AY����ZuL�<�9���W�>A`D�KW�N�4W����u8�zg9h�� Х��?ƷDG�j6Z�������:dxYS�4�����F��,�-gf{�Dg�#2��4�U|�;!\��du�Y:,n
�����|����Yn����֏�K���/�6y�Er.����h%����b>���80�~_3���տ�3��M��[CP�8�2��=��e2dD��:�N����dM$���O|xM�nG�4�Qь�<7�R�7M8R�zR��u�33�ĳ����r���4��״<�^���㲢J�
<&�'r������\��h��&��ʡ������Ҁ*�M�EN<�|�.�] �fr��r֓Kֱ��+W*SI����c{��[>���;�ӺqRų{nP0�Q�:���(@ǎW�9!�h!�w�#b�`:�L�C��Ng�Z�0�G6Uq�]N4C�i"V�g$5�{0-����k��cГȓ,p�����u8�gl�o���a�A�	�������O�Z5JJ�]�1m���Ӻ_-�4��[W�-OI�\y��{����]�����6���OJ�+�Oq+�:�,�!����-cl�$��a�����	�� ������y�(�+���Ȟ Jd�6���!8K�Q���7T"i��k��X�w9��E�q|�p��R���~i~ة+i*9R=9����˖p9^��2�H M
gG�+�S:��s���b��~�~W,�V[df��������$+\g|�'H<��\�ـtoy����Y��'�ł�.ju*��ס�q�ŊIg���%�ɖM���X<�u[0�̀��t�B��vth=|Y�ä�;{��N�y@M�~�L�D�X�a31>���ҽ})_���.�����{^�Eܧ!�Sf%(짱��*����b�8p���! �tX�Rœ��1� �i���3��g�v�W�a���c��M��J���T�/���>�'A|��bS��ͮB���$o����l�C�4d[3���H\hyT��~I�$U���]��ct��N�5p������\SX4���r��ު�sp�d�yF�؉|>����W�����S1����^vq���MWp��,�o�t��5���4ef��_ߝ�_g��_t��wV�Ԙ�`������
jX��g@�,��\5Y9�'��|a� Nf�� ����C?������5�z�-��R�nۇ�Hik� Q�s�.�b��p��G�Be#���Ya���D3�KU���+��A˝�����7�6���\S�Lso�(d��d�Es�`��#�F��4r#�c����t�/p6��(���N��w~�W/�D�j#�
�:��7 �3��3�X}�����j�����O0��j���q̏:������	�֭�O�S��>�5�h�S!�x���D��u�;�&in��E����-y�
/mX#�>Z?WM�7���3�b��b�@/=�{�(��@7�m�I۾)K	T`{�꿒�����M;�f�����3�U�G���^F���͔��'����zȉ�0�Ǯ����G������*/"|�����̦�	���l��Du�Ḳ��Y��y,-�i��^=HK�lerxMk��a�S��j�#�_7N�n�HVn\)���,+D�R[�o�|��kjB�7T��dWZ��Ȩ7�kD�ݘ��7O�7傐�3f5G�,�Jy����z-x?oK�e��^0�7���6I3�q�Jl/vZ*nl�侖���0!�#E�`h��C�m�[T�bo��"���ƌ韵f^Ƹ���PT�cQ�����H�%~��ȕGtj�}�$��MN�?Q�ʳ>Db�:;�X��3�Юx�R;3�B�  ��`��WkWO�G���Q�GZ��{���:1�E��51���%lƗX��KVS
{���'�v�|NA�yJ׆�C`9��Na��B��HS)�ِ�Y�X~��:i��H~Ow?A}Dx�JO����6X��Û�F���);�XW�­"���e1�_�x��em# 90��W.-E�!�O��.�GS,jBg����)Eq�\��XE��$v��6����CZ^ȟe�3��n�r��:�Z�	&��;3�n���Jʬ3 \�X��x��� ��7_4��wJV6nv%ˠ�7�@�I���x�x�n��5�D՞B��0��1J�<�P��1w#�8TZ�p�����;E7Eo�Z�cP$Ch;0��tFK�*[(�؟�^����@o&���	bj��#U)eKcL�(|��I^��BP��)��$��*m����,�;g���Տ1;�h����1Tl���;-���#M���W�VL�2�YF��It1$�ݺr��l|T���K�'Mx�V��)���s�H;G��)�fU���zrH�5�&Z/�A
&����KX�wH����<y�#,_����5����7��ۢ�)bc�!�'b���u镵ۍ��L!� ��u1b�e~�Oq�h?@(��М͗���Q���S7m��1ȜL�}Y(A��1l�zQ?��x��!������ڑ�N��z��۬��9�@�	N��Ŏ��*8�q�ϛ�B���wf#u�W��YǍѠ�v_;&g^��L�Q��j֕�N�}���ǚ�i�%�PH�1�_k�����p)4�,��� �8Y��r�|e���m���M�u����.���Kyϸ�ʟ��=(p��;����\	�9,� U�h^�S���3�R�-�Dn��#�x��۫���[��{t_	�O0�B�F� �y��H[�J5&����7��a{f�-��|���ޝ"`pz��ک".U>X]Pt׉N��ճۏ�W�R�P&+��9�{��&�u� 4�f�v�>�	-�Ed�?	����@Ѿ�}Jp�`�Fo6B��KW��TKu�����a"�9�C�z����Q[o���r�C�X_Sq�������K/��"�$��y�}���9{ln��M�z{Y
�*"/W!��(��{M����i�!�)(}��Xה�C}܇�����t2>���Z.=�
	�}/ ��Π���H��=����V���C��zc�R��#�K�]/6?,�U���L�a��ppB�M�ܓ JI(-ɦjT����@lO�)Ҭ�p�q��`}5}�����a���CSQG��]�]�d�	��z�X���Ib[
ic�=�"��� 	����cI��k�4���^����/�����#����BC�-��U�=����	B��Qm�3~g�Y+��q'����%�#��[�T���Ň�r \M��U�ey?�ZA��i�0�d����u-H��G�xn���^�٤�g1���L��*{p�>J�V �bs��[�ƶ�#��:e;C�m��F�ɟ��k`���(^�j�9i�z��i��kjƽZ���,�>��D�i�S��.j[k`T *⪫��R���s:�dʂxӉD�z���iaG[ܓ��|�s�f.�}��N\8E�0	'���j�c{U�
P��1�Nb~[�C�vq.<-�ӂ�Y��0�}�&+��V��҂lT��+4�/����~��� ���*r��w����J��Z�������������p @t�'�K�)�n@AB$��ev�L{��S2w��:Xi�D�1z�z�������TCDN_a��\����'��/���f%�Q�X� �gңH��ea�"���y�!�1�Nѷ@�]߅������+=�<#�������"��^�UA�4�����&��^T��fm�3�@����S�q��L�B$�݃��O��$��@�?��l,�]n{;�a�����﷘�w���j�%�g׳nB��'?�d���Ԣ��aP��"_b�|a͢L�����#�.?j�͐JB�#YT���p��,��,h�ȥl��bɧ;;¢�G�<���V6�&�\�,`Ly�*�<����O Rks��@ aw�\NM-��=��X�_��~^�Yc�8=@�ߘ�H�ǈ��#}�7iL�l9��Fx�V�5����DK_n�&����	)�c�$Dil6��v��/q��"��N��P:�RpP�,�"%C{�ԭ�:�/o��02��� �<��B8�{$������o�7{��§A��V3�Y�|�L�-3�p&#���Q���	c	����j�XH%a�􊱏���nJ�vnX&�W��>z�|V��F=������鉽FJ�Y;PW�R|�8���|3�Iٞ��r��p���X/9A*$@�B�O���%�|V�"�?�L_��
c2r_��� Թ�Zr��!��Gr�6Di��,j=!�:�>��0�U>++�N���Ǣ��}=�;��;�+-/ů�I`����Pb���q/�meY�eںl;K�Ll&�Į�gD`����;�_�/�2Xb�w��Ђ��������j?h�X��y���n�h���)����Ԯ� M��8��:��@ �L��������]��t������ S�a"QY���l ���M�O	�����҅>�[���g����؏	���¦����t8��MΎ�z~jM�M�زo���Wv⃫Kr���?�4l	L�A�=�����l/*�\5�Nʤv=T�j;'�T��B���׻�k���]����p}V��MZ��qB��FC���u�9�^8	�t��Y1C�C�8Lvo�Q���T$ߑmd��&w�1�AM~F`�׮��( {��Η�J��-���d�(��؛�K�D���[��}l��)�mz���-�g�_Z���(A���u�gJ��.5�LC��g0�'\0���"V2G��W�>2�X����f�y�^DNe�w�"�(Y��PϿ �ږS7ť8TUt�t�B��m�O��D��s'�(�P���C:�G�����x]����Kj�_u�����}��h�rd	%>#>�1��:�
N9au�0�ͬ@t82釺A�O��"��фo�?�1Y�$�<!c���'�*)Q7D��S�����Ƕ��U�<u7��Ҋ�
�#�i����+�����Q�'���H�|������5�4#?��kn��o�Y��ň���H��L�A�mM������tP�7i���#�O�7�qƑ߁�2XE_�F��{��JM2Q��ܵR���G��sL׿��֤���%�H�n�f��􀑍�@��d��������p�S�h7L��9笨ԯ��jߢ��[������5e���B�֠�����Mڲu�E����dRn<����&�̙N�,�7܆�K��r�#�j������Z�B��f�p�?	��;�l"�%�7�����R����F���G���ܒ�|������P�:�5o�'͵U�Y28���-M|$����L�pȹ��Q���O߄��|~ѝp.?�*�D=��R����42����7UΊ7&�� n_��珠��:y��{�2��R�	���ؗI�Q0hB�Tm�+�I��������~{<�����D���^P��֋`���m��&�c�s6��ۛ����N9�s��:�mdL$�]7������&��b�F��bR�GN�$�I�uj�&��}�Xdw���4¶�>��k9x�8���^���K��w=��dc4x�Ú�R��ή�# ��#�hg��f�h����$�$�-vހ�{�
>/�Q����շ F�]�"��8�-�0n�O��|��7��1��SM�Y9�ҳ�bi���Æ�,�p%
��v��Yn��M$��:ͱ`Y�2�A�Aa�p*�AG��,��c���5��Ew!T�Q�Dp_�D�\�%Q��Z@C�RkD�5�峉Fp(�����l7N���n3O�X߽�@��:��r�=�-�A�d��?M}��G.[�R�q�Fo,�gT�wenuj�����e�t�ǖ=rG��v1�/�)U
� ��}0�48x�\{�4�u����p:�%�W,�B�!<���;��O�~)j��*�F�s�2X�VEb̃P���y9q7=�+y:��C�1֌�r#m?�9տ����a��4p�6}=�0݌[	^H�ľ��x���..��в"w�p,�X����`�K�{�U�a��m�������z������o�+ |lř����.C����!̑�L��r�[��@�'�s��B"��:Q�`l6���x�!�
��m��N���#�z%v-�i�X
 �*JȨK	�2]��aog:�%�:��	~cI��G���A��_80[$Qu[�|�1}��f��u/���%�nq��i��i���O���h���ӗ������Z]��K�C���a�<��`s�v[�{x��oS�Y[yV��&L5rh�>�����M@�Z���.�;4ҁ5G��R�p��#���J�T�5��4f�$pj����.�-���rI<J	�QIH0������⌊ysgdw�q�o�	@i�su��]���'��bK؉Pv�N˙�X����pm1�(����y����26�k��w��5%R8���~�d�1E�xk�yC$4O�ɿl��Q�]�W]��m]��J�j�S���:����g�yR�hJ���YE�S���G����}�O�G�:(�V��Qz�o���E^~��`w�r��I�DB�E����-j=lq����F��C�+�n��M��̼K�["�#�uuI�wV�'�]�l����U���"1g����,@��<W\���v��>\%�T��&��Rr���!���J��=��t��lB��aT|�.ev��u@Q�<�%&L:��C�p+�1�:�\�u������G� �b�N1�P^`��,��Id~�۬�M?�A���*p�r8Y�HV���b���3GD�(��A�څ�R;��db� ���v��<�8����r$�lcHP�����GY��eP�]�[�,��)Z��*����G��H�+��0i�^�u�8.��.��H�n�i+��k�W���R%�X���,����QR�3�-
V2x���B�3�j��e�dl��خp^�ؕ\8�͘�M8�ڞ43�݁�{C���F0��g['��=|�ˏm����̭F%�<��VMi;��ܴ/��?ٷ�(��Q/�ڨ,/��'nY��}S����A��r����5��T�ڸ�f;vc����k����c0ex5@ ���1��A��N���+�-a��74A�����w�gGR��m���wP=�r���*yߜ1�p �W��5��(��tg�N��f�,����5"�TߑT"C�e!J�&n�o�	2��1�;�8�7����َȸ>�4JWu�+��a9�*�(�!Y_9m@�����%��;UY�br�O��M��`6��a	�=��1K�!�œVf��>y�z3p�BD�);�K���D��2���xɽ%��?��4��J^�Rb���#}QGB������+"h"�Lr��frZ��RQ�,Ei5�"J�
��Ie�s�U��6ƛ��<�MX�!Sߛ�r�;���˅�4mbAp_���.e��.RےY��������" ��l�O�~��#�>� �Ѧt��I\�%����x��vXf25hPSn�I�ݪ�Y�vC��6��Egu,�KAA	�)�SF�n������0�]p�U� PbY4���E����Qg�V����ҳ��{5�%zL
�6O�d�L
R���+<���(�?�R��32�����kV�$c��r���Hb��$�d��Q�)�FT5�hֳ�*���^;��\�h��Jsyt@k�[�����Z
U��*+�J�?��7ږ����HDR����}P���^󹸷�>s��p����?-�\�ڡ���1� fuJ��i���|�w��'jkK�C;�H[���a��IH��2��rs;��m�#%���(���j,āh(N]�bԷn��&w���,����λO&�����6:��ڎ(��oϠ�e�L>H}��3۶�s�K;V�/ɗF�� C�.[��P({��~IA�|6J���a�曧i�&J��;z�u�6m��KZ)�ζ��8h*?���h֌>��{�<l�޽�:J�4r��վc��կ�l��f�Lom��8&�\���d�`��}C3C�]�Z����0�i��u,�i#�n�eݧ��@zJ��%��l�jY�0��)@G�� \�����S�wr_��rԦ:6����ʮ���-Rnt`&���ڎ�7��a��R�w��fK��R���M2���K�ܩ�H��6�G���y���J�sz�8�9Qb��u�:����k\=UJS���ܼn�����ˬ�s��Ɇ)K�IG�[>'|k��b�B��'R���yi�9��u&i���U���9MO��N�e)��=�[3t��}�h�J�sKǄr���[<��n-W��=؜y�i�{���#�j�PA��9t����ŗ%���E!��ǧ&
���We�[lm��uh�\��b�F^����@�҈6�\�0OGb�7?F�K1:+����aɖ�S�/�D�gLe�p�/��������Rm�f�,y�:x\��-��4�9���.��m��-=�0��k6�e;IҘ$�v�x�.ׂ����I4u��cxцb4�I�(N?�dOܙZ��w)ίU9%#܇';p���{r�,�vYR���+���:��4h��ܿ;�d�7J���d~�S�I��Z�Ȉ�9S�A�p����ߚ���nӳ���J $ϑ ��i���D�Жɖ��'�-���Q~��H?���A&�JqBLȯ��zKQ��t�sp���f���Z�"��t?2�4�;Ɔ)�c��/�5��)AeWc8������&��~rWj]I��΁'4i��;,1�_4�ޙ3��Q�d����O�9R�;n���Ņ����>��!u.c�J� ����_ҧ�ն������W10���}�^�}_�O�F�)�5�>�����V-"-m\�Ҧ��ߥPJ_��� ��횧�6%��-p[��ׄ!���qH�?��~L]�s�r4���".��3��o7�@�s;5��m��d��ږ�-�-�r��TC}2L����f��It3N�Hey:�6�[��jt�ԉ�G�������4i\[��2HW�""f�r������_t� M������_Z)~�p������ Cɍ�-�,Ѣާ����,�հ�R��En�kq<*��l��r0J��k'ж{�U��1����R+Z&�B|�ñbݍD��SJ����߷�]�P�K�l�A 2�A���]�|m:7K���Jc�	�[a�y�=ܗ�O�+ͻ^ʀO��%	g4;MNf~�桻1)15�I�~B&$��7vY��xK�SR��7cM��T����\�O�1�oq�$'�M?��;�a&�Dվ^-O6�{����7����jFi�Lj�c�oУ��8��R��&bH'; +A��
���\���a*�X�p��f��&��2%�/�§c~Ɯ!�i�e)�xX6y�Ǫr7���'i�~�j~\�QΕӻp���F��$��$؄���;=A"ۻ�j�s�[�O���/��@I �E�M[r@v�)�Cm{�G�O �?�2Ųi�!���ul0�-�2�aA"/:G��.Q�N #�36D.�b��#���R���,@�Kg�و�߰���P'�I4�lF�r�٩�0�����廬Or�R�qϢ�����>��<F�l�e {���=$�09�Dau���� �d�&:���"�}Qn�k�>0ZU��]�ZfW�(te��\K7�����9F��>���`s�
�5�H!` �N)��1?��kd�f8x���HA�5�����-�J��خ�"�Ddt9��C��Vi
Vj����H�*M"���x�dJ��T�R_"t���$g�h�7�f������	!������.-�*]UZF�X��Q\)��&%E19`��(`�^���s�_���ף�K��#����R�c?�_np%LV��n���3*�X�쵸b4����E��k�'Z@@
�p��.��$�f�OԌ��3a����UD)�Gɟ�A`DH���to��b����jp�w���nI�^�ݙ�k�9����(c��ܞj"Y�)������h�]
[+�s��rY��X��Oԑ,�R
5zRs��|�0��8w�oO"?�Us�~��!��68aQc�������M���[����;�r��
ǀ�c��	Z�$ iP��Ŝ�Y��j�:���Ѡ���/�f"5Z��%��	�ʠo[B�`�E��Y����r��j�=^$1�^�9x�7L��ZՀ%���mܭw{;��w�GzO���n=�7z�Z�%5�;Q�gQ�Ӂ��5�E����M��0Ҕ������i�\�ZsV=�&��� ��v��	�/A&w	�R�-}{��/"�Ms`&&�]Rl��n�x�N8�_�㮼���DE����yw��d��y��!
��]7* f������J�I3����>9��x#EU���(�-�Ba��K�$���rʮʺqPp�'"���J�G_�,�-WVf:,����"W<Y�����{@ �V�U���$�Q��$���ƞǚ�t�SfJh�$@��k�n�]u�w���YR5��+<� 7�Ϥb"����� \z(�/l?ߠ����!�g��q+v&@ �k��g��y���6�����u5<�s�$�����m�i<,�G3�m[O�*�Xĩ�k;r	\�#8�oQ���69Te|� f�U羋:�$,*v�+����c�t��V�~h^�1�&;�bC�=whe�$r*4ьf��S-ˮU�	�So������P�[�g;Jg��-���E���X�V�}l�'�@��d�X�َ�Q ��?3�K��
n#88�-q���k�28t $%����6��:�H�u��{J8=�Mc�G�Jeo.M".(1Y���t�|�٥��I��h��B�TL���D�6X�Z`��?�.�ރ�Ay��s�0]�Q_�F�����t��ER�w:�xE b��<�2��� �YrD�܎\�#���;�%5�ª?�`�ܗ�Jj�&5��';�JfӤ�%��.�GsZ(�%0�e���0�	'a��ٞ�@��Q����K<��{���A�lr\�LK�0�c��)����^��[ȃN^���4*�Jƙ�TB6q��H���0���Kl�K�#�m���Ma���n��M�Ɖ����_��E���X�U����'D�p}Z-�y�B�4qҺ+Pq�� Zp�CCB��0R����$U�}R�e�kt�'��J!�H���>�_���"�*U9�{�.��Y�<:BЄN���>�.Ut�������x1R�<��
P5���K����� ��>3���c�xqqN�&	�`dd����`�Sм���w�:#$��e�F�*0e���?�@C�ա�n�JGn����gKU���	�2�(��M)P�v�YŮ���1���a�q>�Y�۠B	W��w����3s�1@	[v�0G7t� N�H1Yc�,��V�J�k�y,�b����Z���5!�в���9�J+��96<ӝm�F�z�W�у�����.ƒ� �U듩��]7�h�ԃm�5d�� ?���ڔ���5%�V��㣄{��$H�lY�І۪����z��g%�����Y�6�T���;�aK3[������\���L\�a��U��`�����W��G[�8�D's��S�f�W��s�����2�j8.gF�˫�M�VGU\-��u�o�_a����F���dnFÂ7��s���	Ә�;V���N���t;O��P_zE�<<Q�����90�-���o��:�	PC���M�a%ڤ��@;9#�
��z��ԋĠ�`KF���Q��<�?�e���>(!v��ڷ�����:΃��2���]MW�|��_yZ� \�T�d#�`[ʋ>MW�'�)�']��ܡ��D.�&� 8��� 8�&%m�'+�M|��^f;�T��/���c�����?�@�<�5�!1Dh��u(<ډI"/�5�`&3�l�p�
�jf�sV@�8ߓ)p�9j�B��/X�sO�g�e��~&DJK��Pؽ �k�Kd1<g��y�"�T~N1 ��b���Q ���:e++Z��%��v�ŕ��F��t��ӹ�\���jY�EO�7�0�j� 
��G��٢�
���M�(>�.�~G�N���-wf�S�Z�Uu�|�1.�6�"q
h��q�6 �ʘ���P�M�����dC�?���T?��y
���i�6&���K�]��'R���66����K].f�P���Oo�t������^:0�h�/*���(�����M<��a��m������$�6��vx�O�U=b�k����pO 3#��z��h���j��EG�E3���q�v#r&ĖOJq��Tǋ��)����k#�#�#><�W���]�~��1o2���a��z���ӌ�&��h?^�,��qZ�$r�p��qsx���x��a�
T�,6��������6�^�� �-�Y�vM�I-D<v٪�����۸�/��WV\�٬dky.�>��xߎj�c�րO�F�)�4|&�+���5h��-x�;:�"Q���K��m��7�c�Qbǁ��rׅ;b)ꊁN�BS��Ը�mjZp�k�.98|��g�N�t���P�e��^!���X�pM��^j|��BN%��1��*Hp�=��C�qdsa����u0�+` :�w�-}�*��m겷�B��}�
PW	c�����\�^eO3[���!Q_�*����̀��hw��=�
����bx����1w^��v�CO@��.���̙�hA�Ϥ5r\�����#��-GǨF���=�3�����b3��� �_�?�ʋH�B��!6��fb��n.\�D`չ��x�5�E&;$�bp��iaP��춏�1��P%�%�7��*\�LcMNmP�u�Fm=9L˂LW�u���.�_uO�A[}6?ǡ�J9�Ը�,z�RdW8��XnG��_�C�=C��u��6n9�Ћt�J�c{�v���x_)���s��%ـ��-�Un�5�,���47P�yk���%:+}'�=���$�ę�CG�h9Ү�*w��V�T���e�;K��������E��Z�hBXf�0H6 ���I��P�9��g�Z�2�D�%�@{�8K�:I��}o6A��Ad�6�{�;��܅E��T����QݳMƹ�w�T�ےuud�V��H͔JmQܼ���W���%s���Z�EN$�5�sEc9̜����˱�X���4!�� �7�e�1���4��M(�8nH֏T�n����eV�~�a�� ���DӺ���î�����΀4����
~� #'��d�-�	=�ln��q�#ᓊ�̲��P+ �\���7�ss�yG����M�\{���~�� �A Ră� Z}wh�.r��vX5�"�Q�7��e��_ʙy��G΂��Ņ�Z	#�"���?Q("cbQ�$�0�֤�b���6���T�RCz��*��I,���,��?"@�}��QϹ���k�g�	WB��4IR{��b�4��y<����_R����:���|��πQ3�\��%*��o=,�m����ꎁ�-*P�+� ��*�\I���O�br�Q�-.5���,go2��|<:��t�g� ��T/�(�\\�	���t�I)��*���M-��w��xG|�d�=ݫ�v��¤���>��05���iɧ�ٶa�����n�l��6xoj2������$�	n��Jh�9�?�q����?jC�{u�k���c"�� $Ë��ʅ f�{�g���cW�ikf��%�0R���¨@�K+ � s>���4�C�N5Xr듩���Y����z�
b�^��m���ή�{I m8���Ha��%���û���OG���w�鶒O!@�o��V!��A~�k�J��h�/�d��\��5���W3��1�}�?W���
���%U�Gq8��z˙�����ryu�ǒ���u���7`�*�Ք�>�j���/MJ��n3��q {.d�U"J��k�S�G]��B��	�"/�a=f8�Ph�1D�k-�<	�_����m���$^rE�����8�{�B�ZJE�Њ㓝�R�\c�ic����E����`O��T��>sMp�zRk؞C�k��<P	�&h�B e������>'��u���ǁ�Q��XN���ق�*� ?�:�	�
hy�2mM8=��R&�W���]�٠g:�Fh�#�v� KU�E/���9���(D�6�Z�'��3�S`�<j�lZ;0���V�hsD	p�(Bӄ��K�׿\K׃�H����S�������W����2O���0�g����X݌�v2�/� LE{?-t�ҍg���{�FN�j����K�!C���L�գ @.�Ē��<V �|�g
	t(��y�Moz!	�e;�<�~Y�}լ�)�&>��4�e�M̈�W�2z��{�(wΛ��*�m�!���\�j��L�[1t�&�>I�?N�՞l���������!�8�`��	a[��:8�"^���.W��i��_�r%�t\�7J�߷?�v?����f�b�ǆ�xv�U�
���:�LN�p�?�դ�:�O�!�����4��.^��=)��{> Um M�I�".�-�5����(�9c��^����G�(G;�05�]qZӣ/��{{�l}"A)D�Ҷ3�eL�(e;�WIW�����)�;�����mhWI\�9�H���/��B��UU�Q�֮G�(.�)J�'H�6V����0�7�yy!s�&�wU0�Y��V��_�Q�F璶��_�6��EzHXĪ���"���m��9t[�X1�/�OT�	|Q;ۦ�4��	|*��j�x�#-�!�\�<:˾٫�1���'Cޟ�n �#z�ҫT�Ԓ�����"S�����ZЇ !��fa�4�F��B` �;��(�4��3WOV2��M���0@�;��zōuԡ���u��y��d�o����◽�P����� \���qpH��V<.A\�q�0J�+�AH�K�5T�0L[��T�p�:������ �a�CP4�߮��3*]OF�#�������G �%�Bt&�ck��@��ǫ
���ٯ9�jskwK6�%�S���o>ݽ湵i��`Jd=|���Gq��Xs�GZ��C��xX
�*��E���y�Cq��p���C��Վ�Xa���p������cYP9z;��g�ϯ5�gi9�j��'V�:yg��a��B@�ƧV�08��,iF@���&4��a1bR#'�����FG*BTgZB����Եi��E5˴=���-N��y��?^����Ţ/����oH�"+jQ��
�������D�? 6��b3����i�ǻ&Ly�,�Qǁo?Ɵ��Ի@;7Łn�L������~捻�|Ye`�8�T��4R�FL��fZ|C�P|�ѝ7{d��ٜO�5_9�=(6Q�.���'}F~�����I���"~�K�5�oW~* ��CN�¯o]�B�+4_Eu�.g�Ʃ����b�����l )�	�k��\Ǥ�7�U}um��MI��s��{.��]<X:�ީ�N���_�+g�����@li1Ya	Ag���u�L	�J�X�`?3���ݗ}׵5���N��Ue���J?�O���yw}��u�%�"櫶KLX-��=ءRHA�n�e�;�FA�{��iK3�I%��T��r��UF΁�j�8�"O���܅/'�ehؚ�d�GlfUݼIvcL�E�����0E��5������ 9�{rK��f�/�x�{�Z��,���lA��xf��㸵�YN��@�D��]&�l�z?#Ĺ�K'z��:	"&��1W�)��!SN^��Mp��?��\[�N�0�&�*)�R&���p���|qV���eQ]��/�毺@Ll!�@���x#���b莞�*m2},��ۅ�7�?���	�p��+�8=n���3Q�@��,�87 �D�x8ڥQV�y�0�DZϜ���T���Bv��������$<c��v2�%�f�ԶȦ?t��d�ϱ&P��R%��IZ�$�c�܅�չ"��:�yY�D��X+���d��F�~�JeN�������wW��w�ԅ���l�^Q6Ni�cv��G{9����=<�&g�>Z� ,�q�IhL����ƫ�{!�ok˹V73�:��W���	�{�GR��e�]�x?�wv�TYY)s�Mw�ڣ{��hG�@��>$Ʃ~z��6��������s"����t��Fz�KW���A����/HM��Ģy<��F.'�	���熙�	���T���kq�x5E��'里�P�0`�g�ЦEf�4�s���`�P�B�����E���t����&��KOm�s��rG?}�7y��[��>`�r���₫K�h������G3��|J0�II�p2E/ڢ���g�@���T����g��<wae��k8q�d� 2���[A�t�Ũ�Pa�De���T��&i�z�D`�!�,+�<��_�$?�%t�a!�½�Z��S-!�b��A'��A�UR[q��u�׍T�T��pJ��72��%��S�ы�|Կ�5j7Rؗq[�� Kb���v]�Z�,q���N@v���o�X0؄���-i��Xu¯���Y�H��NrH+����^�t�HȜŚ����<�vk��wRg&���."ȹ+q汩ϻa�A�A8������/�-7�Xp��y��:sw���ǔ�����}`S5!?��_����o^�k�\�M�;{j��w��S{)�k���O����?�?Nf��$�s�S���P��ۗ�Bb�Hݔ�;�j�58�Rm�x� E��x�0�Jc����A���(w�#�SF	D�G�k�K�SZ��3S�a?�'���8��,C[�����DK~ ������<�m�#Kt�������2&�Ϣ��<:E��؟��Xػ��[�]�߇��76BOqF���F�P�BR�e^���{���\��{��u*Ut���?�_>47��U�J�������gͳq	�����D�٤�;'�2B����o����_2�bw��;R#g�vFֽQ�y���fJJ�vc�^6 �T'e�;=�Ad��ju%�	��pi��yÀ��8� &��vD,P*�4�ρG�ނ8��}gB��d�v~�B(���}A�tdE�h�$�iU�ك�4.Bm+Qz5̗�Z�+�Һ4�,/��ZzgLaLx�H/�P#e���$��,P�T�>&a���*8�Z�D0&�Y3e�`e"!ԑ��E(�
u؀V��@�ΰql��N���ZR����)Py6�j&�:�8�O1.�3��y����r>x��K��$����*��c�H�ݢ�-��A�g>�ˆ=��! �K(/{$�?��3D��IE�$�Z4\���H�Ү��^H&?�8�[wkU+���ޱ��tQ��F��sU�M��_��5����p|Dc�[�z�M�^Q��F=�]K��i��af��M��_�NT����禀��s���7�?��7��6�~k'<Nz�n:�HQ�6�����M%w��Q�b`��3?X��!�{5)���X������E/5���7A.�j��`��*�B��1V��g�#�9�F�Q��Shb�ȩg'4qP��3�hQ��i�w	{n!�OfX��m�0n65t�-:أQx0��Kz���
8�{���k����	E�(�Yq��[82 �9z�ɼ�p�p�eB�,-�!��n��o"��%w�u�`�l�B5.��"	�����~�:3�3Dԛ���
�l��S�w{``�O���+u���Я���1��j��o��?X�DC㺹.A��
�Hj��[�5E�)���Of���,�Zp��-�犅���p����;�wĔ��h}�̕N�"�N�L<���?����Ȱ���[Q]d���]�NH�W�s噚�S�Um�����t����qT\Ny��Q��=�]p �d$�|�*���wl�{��KR�E�lۋ�I �/ՁЈmS,�Ns B��g���߁�\�j�Eb�K��Bs����G)^�D5ɌM�w����0𻀩9~h4��8�N��U���9 ��ѿ��S��� �cw�����x�\�N�r��)�����ښ)��Q��5LJ�(߮$���dL���抣'�y�\;�lj��EV]�sR�P&�x�0��bӅܮ�����8��$F�A�gB�P�B�rh����_���WȜ�y��!�Ly�nQ��U��\Rr.v1��G�W�ԋTQ�7��.h��C��~Y�UUAo����elo� x��y�yq=֚~In��R��G-��{�����v����aXT���Pao���9>�(#�-�(n�sM��J�I�Ά�l�N��{r�Q�ފ�gk�@���&�&1�-�A5��5� ��,�3^I\&�?:��;��zg+!�^ܳ��"RU4Z7�<�ՠ��i`���tN�?��:���Ȕl9E��	��4�]2^LN$
�wc�ϱ��〺\�\L'�^yfjr��]����c�ꑜ�q����k�W���'�ǲ��p�K�c%;��c\�N3λ�d��C겡���B�c�h���Y�vy3����:B̎���ݻ�-v��Q�z�,��[:Bd�Gy�/�;c6�Ǌ�A�{CS�6H �<E�ڠ&ҽT�����B����)����}5�H�	J׻O-/�Q]Qnp��+G������/�[��>�h��-]�+��@�ٍ����8���]�7�>1j|�},XM��eks���;@�,��5a�[;s�uhJ0_����t���Wk�"�u�����J�s"L2z���ij��9���(w�4��L�4:��sEA� �?�t~1��f��b���.��ť���;��σྀ��]GZ�T '�PUl�L1�?y��'�W����g{���1G�n��=[jڏ���+��
c�κ�z��{	����p��\�%���B
	v��=#�E�D��va�t �d}�0h<��[â�"}}��� � ����)R�Eq�'4P�+�Z\)�I�.�bB�S���W�l��G ��o?�ǧj_<�i;��b5�
�?ǊcQ��ڷ%W�,��`b����S�|B��=F.�ZX}e�$�m��*r�V��;R���l��Z6�a@��e����ҋ4$��%�P
���8R&w�W�\fc�����:9WB	�m��i�7xV����;�/��+�x��@.����}�2��W��O�U{) s�E\��q!q�A\��5uJ��5� ;�����o!�S'��x�A�1��w��:Bz�wN�:>�E�}�C���!��83@�s׏)d	��6��W�*�iK��?��4X���Y�j���~���h.#AL�p������9νd}��Hs6�F$���/�����!�y�ʿ2.���&jc9�T�C  ��!x�`�sX�4'����y	mjޜ5��*[U:iA}d V�t-�U�Q��>��B�+�@����hԲـ�.�8����-;:�n^�r#/��.<��o�����
��b#G��Կ��H�&~3cSjF��M4��E(F��d	`�e��EnC\9z^U�v~֣b)�Da��
u�3������F�g+���.�����ZϠ�y��uL�텗4��m(�������Ynk����<f��^��F���Ŭ0��,���S�'n����⒚����<�ֵ�Bb-���V����)t�����ɹ��0c>H��j:C���C�O�q���;��~�p�?۶ӎ>̃*qR�gռ�tA:cF�O�O�w	�Q�Y{�0�h���� �q�ݿAL�p��i&yt�1�2;Y�3��3Pj�����Т-.d �;�ai48ZC�c���I��@K ����`�� �������q�-�8��ï�.�YX_2�|{��G �)Dfam�T�*�n{�|���i٘%�C�0����q�n�5g=�s�>d��~~M���Ff�

p ��{
��O9�S��I��CJ����>���b~q��$�������U.�E |H���Vtj���Ɨ�4]���8����=��>�3�<6���$!����O�&T�Uםl��vf7��M��i4�Am��'oD�[��y9/D�dԭ`e���-ӆ�;�]z]0͟��uB�z�O��t��f͵Ľ��
�=�'�����G�q�U)-P����ŵ~J6���p~�E�~4����[�� ظ2�@G��3��ﶁ\���.� ���c�)��b�XX�YS3��b�@�����p2����ڼ�hWE���B�Tׇ�s !LĈI;A�@�yk��	��3��Ο�Q�1x�+����L���"K�T'��@33�&�<��{ͩ�y�w���)
����6�;f�Ri/yyU�Y�M7�lc�$)tn�T�|9�����3�w��=�jO u�+��n�5A�+�����RQ�E]�.�{�7�Q<R���LA�S��xۃ��щ)���s:f���8��<�~�	�a�6��F)��9�@PC��v�
ټd�CW#�m�8�?(iv+^���~ęnO�����ln�9o尣������m=8��?��o5����Y�=a��yo]Ơ����h��]w�rH�oK��2y���Of�|���������M������ٰX�o�)G/���"`~$�m��G��	K��ֆ�r	^C�?A4g���#�[*k�퇴(�	i��N�_��`w\��[�G#ϓ�����X�5�&���o<K���K����&�[�i��х7�d�F�h�M��\�t�˄����~��m<e�ƬGTh�����8%^��b@=�����h���/]�D�I�t�.��&�&؋��-�є{\
(�'Ŧ9�,�~���P����)�)���2 �wr��T�m�	�8���s��?i���*J��j�"�]Jp����ӷ��_[����6����"5�#d�/S����a�1�K�9��B�[V�(�y�[�$���e<��8�J����B��6�߶�!� ��V���k�����C��N�B��������vm�}�67[=���F��f�يZ���?ꑇ¹�|��{�ESeX���ғo9����
�e<L-i�qR�8���7�\9X0��pR�i�E�	�'��l�^.��8˕�۩#��,9��DIc?��	�b3���ӊ`���z#X�A1a�lG8Ӑ��I�Gu��q���aT�ߊj�<���k=��*�VT�
�h�Z`��G�QX���Kb��d�A�#�k�w�VZ��=��\rD}�ZI�uc����;���4��IJ�,���$��J���ݠ.�>6j |z���.���VH-�{�X�@��z��$�e������-`n�x��b�R<9P`U�Կ��C���BMO��얌=tzq�I:r�4ݘ�&����C��)d�9�av���y���-��O�{����5�qv��}.d���A�HU�z�	�9x�;P�/gf��]�������? �I�Y�J��й�g1K;��S� ��Ӻh!�L���cH�g8+���sSd
n��Ż�_�=���tp���H�	�*�$*���y�M�7��?V��C#�<�X0������֬�z��t!��$��r&׶�ntP�{>��]p���X%Nm×�D�SE�ϵ�8	9���ī?���\��#`h7���_�.-�7M�$�?��ʊi@���mfJ|��u<���wOtNA�4�F�N���ն�0HG�k�m_���K�W��^	�Zbgf�^4�N�^��e�}K����IOˈ�Nvdi�$������,d�����~JR>�&eraS�N`j���ޙ�A�_Α<���H����)�¤<R{zk~��h�iO@͛ۘz��3�߾#�{G��b�@�VV��[�����# ���B�+H4k�W��K������<ݣ]f)P8iIr]m�-�hD�7-T@�ci��7t�6Q�T�eʰ�CC>I��:�RH�q�)>�AJ(�U}��Z���g�^��Մ��c�u"�A/�`��k�ԁ;J)����h�ڃ]���-�=��\g=p<΋�H�,���a��5�<�!��%���gR��|��ڣ֍t\~�΢�:��x�ߐ���y����9B	�!�ɤ����w��xK���#��c�%2���R����rY;T�	��f���/�n�Ȏܥ^^��B?���#q���Z�\X��Q �OJ��$���brQ;{�S�H^U�0)IU�:[Mx~������3��%j*/m�&!�aM���+���{1�Y6�](��B��%Z�ׇ��^d�wu �%k��8��K !�j�谇T[��eCAi��C�O������Ƶ�I�4/IF�V�
��&餟q�ց{F�C�q��^k��{ͭ]�O�q�4���I�r�� �_�	_�=���ͧ�y�ԏo�V���AK(S.)��R�Lu�v�$%�L.�e(�#����+�r���KZ۸�ŷ,�w9�j5?��kCT�dى�ԏ'����@HпV	�٩H�^-��C:Кgc�f�Zs�*�����m-�d�D�ݿ��Z�2�]+f�j�vS^����Y#� |-. yi8=��q�i1�w����t.[�"�;L����,rS�����	7�"�.1̲� ����R��u�F�͵}�Z�7W��o$m��nːZ�i�O��^=#~��e5d'��~=�Hw�����[(��= -�0�`^���� r��һ��J�?-�a�Ev��u�	�x���fZnJ�n s�#���r (�9��g�9�L�N�h|�N�W��f���
�qդ�q�LH ���7�/;��ܱK�5J��c����@�tK�ۣv����SXr%��9�l�?�E���q(۲�j��E�@���ˇr�*Adqu����v?:���@-0��� wc�<�u�����r#E����	� fu���i3�Exk����丹�I\9c�4�*���F�K�+�\c��	^�z�R�ې�ڌ�=��6��~�/��oi�a�E�1'=�= �j��c�+i���W�Zߕ�V����t3]֢j�å	;����K7�i#&�t��jx�����:�m�T�Wf�����^���I:ES��v�ᬫ_t�Kܹjf�.���vڭtz�Z�E8)A��ӏ>�z9���i�㨑��^ʉ�H5�
{������	O��Wē;=�����1p���g(�I&�b��(&9&MK�&v@�N.�׷幖�@�2�g� 8����Ӊ�m�
����(UH��O}q諘׋��[�����O,p�l�@J��H��X�h�aو����ۨ:կ��:Q�v��7�oA�q�v09����=MTzHN���I���"�~�ƿO@�u>iCF"�z�N��*C���y���8��.�����TBG'ӕK�~z��n�1���\xd���iv�T�ȞÍD���Q���ѧ,F,���;mQ,f���"�f&�� bȆX�P����jP
j�D��)�}��\[$�s�j��	��/x;��ق�q�z��qE�[��ŝ{S�Z�%��e �*��:��C��Hq��-W K��ҪI1ڹrm5�6�}�wr �Lax4�_��zn=�O��L���R�r:!�ުR�?��+˚>>A�u���/�'R��O��lZ�yo����Y�o#� ��JM򭰾�w/�t���
>�����˞�u�%��?)��U�W��_Te^t�&A&��-� ���neJ�����[:����y��51n��^�L�|���Lp���I��X
�=���p^�sE K~�Cٟ�f��:��X�`���\�¸m��3�v�Pz������Xm��� Z�X>;��p%LC�}-Z��v��r��C�H�����?5s^_	�,���9�ft�ha��f7
���F,a�9��b`u�JFgG���@��U��tg��m���pU��D�u�lwcNK�y�0M"7�M�2[(6`;ȏ�3/n����L�L ��D���ˉ&Ϣo�z:Ջ^B�~��%��9o��AXiC�U�����>�����������O.�8��_���f�J�ʈ3�	h�g���T)�V�����9䮋f(��G��b��Zd�7��/$�W`j�{k%�w���(��MC�����_*H�o����Pjc{s=Ug�ڌՙ{�	����@��v-�nF&Hr:�Z|��F��d�6[XI�L_�gΣIy5,�!��Ƶ��4��fn�@�T軌��_�T���l�J�9��HYF�%���m=�! �N��#Ҩ ��#���r��~��U���#�x#�����*E�5���.� ��4ސ�͊��B7�F�&�B�~s�/����u��jPQ�,ū�5P��K.z��'J����,-�u�F�W
�Np���<x5Z(9�H��C�#�ȓ��}�_J�e-��G3#�K�r�<�Ӎ��c.����p5�@<"���aH��t�-ebD �����mW��=Қ��c8D����Cm��יE�I�{c-� }����27/�� �M���(��
�kKΝ�i��C��J<�['z�Gz/���+ ��uSp��o0��4J^Č��c��b=��я��X�C����4�2���Ӎ�4S,��:���6E�J*6���I��
Bt�2���p��I��2����$��o�J @��콼��A�F=��A��5���I��ʈc����j�޻�,j2���嵭%��4�Y'��_����@�����NB�B�[xd�5	����X��и�7ʽ�c��րTA�7��?��/0��0X�*>5�^2ٓ��L����"�4}<�S��d@���$���a�c���gr�1p� �S�HP#�So�R*ۗ�b!|�c����NG�:/�s:�6��q�]�ad��:��[�W�e m8���C�_A�����'�K����O
�#3$���)�z�������oc}9Dƫ��m/|+T�����w�(P`�"?Z+��b!������. �U+?�ϾuW�.��$=�CtX`Mb�B���ƤL4�����!�m��&t괸��ewL�zpáq<����E;i�`U�{ݾ�{M�*F��2V�y$�I#�HǨ9B8&�-���I;���3�2�D!�r0fHg"�&	�a�8��P��>��D~�Y�
i���@Q����j�]�2[���e.=S�3d�w�sи�j�ش0��g���A�ĭ!�{`�$S����J��[WjHee?<��#���,�5��	[`C劀�&R]��wMS:�;Z:��n��)^E�E�Z���/ߎѷUۧlaQ-�%�QPV���W�1�{��ue��'M����d`����ض�p�ԣz����_�z�a�R�v*̤��敽��ڲ�S�J�_*m*6eV�4*Vܤ���k��s;��喊�F���z���I��.f��<�d�����UHpk���p�{P�MymbiM�C��n�:0��|�v���U2/f���UB`�1�c>��X�أ#L����SV�e�2�N��D�Bg�8�4<���dq`��^M3ζ�Vr�f��S���G���T�.�<I0����q D��W���5X�|S�E@�r��d�`
f��7٩�
0-H���V��-85�P3`;0�H:�*���U\(�oL��V+I=��yRQ�C�=��f�L�a2���l�&ٛ\�(�2��{�@Bm{+l�-�u���"�s�Un��B�ߨ��/�b�ϗ��BXBB{�ǈ��3G�lo�"y P�*f1�iB�E
��yE�0+���
A�E^��s�I�0��P)��M-}CB/���SebE55֋�ݳ��#e�)l� R���iZ)�B��N�=����Yi�K��|�����	9<���U��U#��c���� ��<S���d)SĿ�㶜RQi�&��C,����zT����Kth�- 5�t�X3�P?�lJ��tT����B����8��gp�7���&<����,ޛ!쩤�R�;ǐ�����GO3*f��:4%9������ae8�l�Y�%v[�<�*���՜}hy���� N �K����}�1rF��`0gPM�*�5:T�%��Ot��~k�"b�FA4%�K��V8I��=�'���8X�Z% _Ьżd��ks��J������.;W���0�{I/b��ݩ�^�����yb��;^J5�N�X�������^����3_�.8�`�5Bǳuo��E�`IXz~-�v���6Rs#B]A�~���.�}p,dP��Pݴ�*��P�����2\�K]��j��
��۲	������R�q�f�?]�v:ja�M�\�R|R�e�b�����{B���根'�^q͎��5NY�[��F@����jHr6G{����ZE������y���M ��Pv�M0����+����Ŕ��u ��б6u�j��k3�SRF��S���{K��Oh�ǐ��+�A4Z_�_����2�b���)"�W@�DcaN/|��	W�������?�/L�1�����T�����Z�ABi��K�jŋ�A����.�/'�M8D%��)����Ii.���ݘ��J��©١��ɹE��O�������c.޵��9ٕ/K�HB�f	�f&�C��
��'@��}�B��_t�L�
��:�}�� ��!��,F�AQ�\�k���f.����Gc ���`�#e3�Z��,3�5U=�J��	���O����7_!��F��4�D��dn��˂�S���V�\^x���Wr�ro.�c�)�@H�wJ�fRi������S6"F�|P�K�_���u��,95Z�����M�ƥ����@��xQ'h8��h���F�I'��%fJ�������=�)x�!B��{6d���#�ؤ���^x9Co�W�Px��9�P����o�Y���F�S4^�k�/�発s	d�`'X(�MiB�	[HUH�<���A�r�T��r/�TgL%xV5rI��d\�ذ;���Mo�����j�� t���f�uujex��\�ϜM8�\�"
�����v,P"�QV��[���.�ʊ�c�2y-���7���p�:8�����p :�h@��Z̛�^�V�H�z�C�����6q"!L�����3�ipG<Ss�x��w�6�E!���H�I�\NY:��ڈ ��T6�(��YA����/����(�פ�e �22���k x5�ND��]ɮ���4��z��\�m�V�䗉��%M�s�N���a���y�蚨�V��$���=��F�S!M�d�o�IOB�kE�>�.-
�(��&��A')Y��y��R�D+؜�d�M���0}����5�/�������*�����˥���D�E˒3o�+<�w��
"�	l�:�#�� }dǕ�/�7��[��:�c`��o�s����b��Cm���ג��(E��YiD�!��?�8�J�M�Bm�|ђ���<X
o'���d!���I��C�<��zTFʕy�D�b�͊����*C�ۀ{�_#ޭjR�2�rEκ@J� %���B��'��Mh���ud>��Q���G����4�x��[Ǔ���"���C����${ �Dh6�+0ʕ��J���X�x����#�fIf�Hb���<��lke�>{!CS�'��B�� ���ɢ$8d�҅�8@|���{(�G��ӡ+�2g�L~���Øp�k2�$���EK�|u����B�G��-	�e��@���(<����쮅��(qc�v��~�rF��+�
����J0�"7�w7��$<X]�����
��|���筊m��m�ͱ?`Ͳc�%wS(��v�+��?�����@� ����z~JB�ǁ�=�d�ވ����:�;xvr:0��p�6A��,%~��z=\T�*���(uO	xb��ș�"��$X���dM�e��j���*%y�\��������Qރ]׃��V�Q�R]HΖ���6�m0K���rw�|h�0SUv��k�Hy�w�r�����I�a�W0{{���YÄ8���ۨ�(���9u�r�2o,5�����j�˅v���,�c��� �-ʓ6����#FZ/���?^Z%~ڈ��6j�}e\�.6Σ)�(/�Glt���"�?P^�\})m"�� ���ɸ.�4�E�`i�m�۪�K�0�m�R���$f��S��1ϗ��vw��31����\�y*�DHp�2
��/���J����i\��*ʷU7cP?��H4�=�$�8���ϜT&H͍�yOB���=��Ɩ:q.��E��qwC�[��V�wE9��.� C>�1��<�0;)�W[�OҺL�v};�_�G:�1UXo��z�}�^>o�|!���K[�G���!�蟿W ��6uיk�<�0���F������r��k�9]��ȧ���`�kY"��_�!��������P�љ�����zJ��/�hW������ʴ�s' �Cy���C�T#���Z�^�q��2R]���E��#Y�+�����O��M�?4�-�J̽���8f@���������%�(����n�0?��T��o����s.L�-;!Wor+j�@���Zڲ��m𧎺��q���c�~��R5�⸖!�\vh��,���Q�%v	�gh�� � *��ѕ�{�� @�m:^���gVe�4�rve�Z�f�����Nݘ�<lOn���j�,���<��F�m�]�����m����V�
��ᕣ.{�ї�&���OKL[L���\e/�v�0_�[�����Gg��K�:��C�[�c�E#^�ѱ��*�<�qBl �-��
����KSj%�|�#cg�����mS�Sp�M���z�ҕ(e�I��N��-O���q������I}C��xVv��^���)+�Nn�ک��t8���<�$v�(L��'B��w^i��{�Q#��0Tj��z<�����}[	��	�h@�_��H��6��$	�����w���i���3)�o�24ό�e��F�Ⴭ۸+��4_��>ڹ]b��g�V�ӱ+�^�8ڸ�1O{=�e�	a���`רQ�W?�QD�S�s�h��ت ��y��N�翝�k�G��H��C�"8V+�����%NE��{ ��`Ω���[�������KiJ��p~}žS�6�p|�/ĸ@�ޕksp�
SC~66G׋Ò�b��W�[��'m��*��&�h8���Q���X�[�� �
`�[����00#>("�ezvB� T��(�鴗��u����/������j6[�����D�s�r{g�{�� By%QQ�埉�fTBe�1�
%i|����d��ї�#<:�TC����M��1�ɤ'�ؾ<Q0|�
�<R������1s+6���S Ul�� ��/~���)aU�N[�x�z�7Q��%���h%y��+\�X6j���w��V��$�!�㋮79_����|L.��X�Y�I�Ð�ʗ�p��#�_+�Hx^��ء�f)�	��k\dla��һ3�(�޸-����yi�6�����s�h0����/��n��kֺZ��'����e8V|�#��$�4Ǎ1�Q�]�k~�d��4��t�"8n�hXz���xɲ��B�f��O�"�W�:������x%U�w��3_L����yJ�#t�?����PW��n�7.�����m@/>�O�Iq�*��Tn|%��hZ�2w�#hq�� 6��n�`�����r�][o��pZՖ!��Z��� ��C���
߳���-�	�Ϗ���{Ȏ	�v`���3��b֓� LG�Z�E��y�'���[�\���o�� ��2���昌����#����@Q�fV�h ?��җph��<���v�N�I~16	Y�P��0�K`�(o�I��f0�|Z�JLK����0��<�Y�rHST����#O�q�o#�z������U��
�@qǃ�0�奪��Kk��Q����z�W�Y�û���Bnf��+^�-��߅ݕ�Z5�$zKF0�8���l++Є���r]�$�s�d�D�5�����UN���t�φ��n1���!Ռ԰b���2 u^)�s��OS]���Np@��������4���zE=8��6�"'
;�
γuՀ�[ɼ�\YܠJ.���'�)��oyS�n�>�%�\��K����Ů�m9eK�ǚ]���ރ?6/�_"f�<�	7���oW,a���WM��T-t=�����vj�
�u��#�
��$�	�j�7ӌѦ�죴܈�ROY&wP.��7l3�.���TcA��0)�o5�+h�R��v�YiRJ85d_�z���?d�����ϭ��N�A[�-��m'!��*��}?�6E��M��OOV.���,���MYR��h��q�#��� ,>�}Jodz=�(+������,y��4�X�d�|+�O����/�n�YHU~��/ �~.i�sk��
/}��ĕ�G���H[�0c`;���rP��	
%>C��3""���Rȉ�#|q�-��t0f�ז�x-#wO��z(����0��ȶ�-���r���/���CP=h��@�d'�P��	>��[Μ���r��������q~3Lv��ֶ���6 F���H����v0_�SMf2�T����c���ě����� ��e%�6�� *>��k���"��l�Z~�B�C�4_�ܔsd(�?#W��Bf��Jw� ���8X���:cP��ݗL���LY�k	h�LZ�yJ������S���z+�� Yu),oci w��-�)�}��#�93���H�QL��Lw)v�y"j�Q~`䂅_a��o�$���BgT�M@�9�ߩ��23��.ѽ.���B�&�W1��� r[2yeD�֌���)��^1٧�UB+&������)�{$��4+C8�\:_��~���i�b=�_ Gp����jV�,����v�M�U�Y�L��m*U���\�,���
eA�o�o#������"	���#�ܿ����w���tH�z��M �@���W�@�3�d)7Ɂ���(i�9�˓힤(� ��X�4�NVT��J7���p���|�_\s���q�t�����*21Ũ��<���\�(�lL�߹i�GP���a��
i=�xi�K�ӷ8��|)֬ML��i؁����E{�%�\�8�KCv��y��#%٨�T�4T��A>K����,�2#وZ���bo9���Ҋĳ%�Ld�GV����}��%��� Ǫw�80>p� *��T�S�zC?@�d�{v�5ѲG�����k�e�Գk��
��O�;Fc ����$��3�P�u������?��<�H
�\x��>j����'D��֎渘���0�sُ�S���Yx
��5�����,q�)�`_�P�5��h)��Ѧ�����:-�������gr�,�$�P�F�M�8�T�ꈺ�<05�@�e>wX�S����8��?�L��VQ���-�I�"�-|pL�x�2��$s�����g6b��1�K��L��ө�6uV�Y	�σ]6��%l�����h�ب�7����=��_.��VS��/��ă��f޺��˕|�b G��y'��<"�l�!���*�9p�S�	>�颕�x��1BN�����^�/��t5��*�����A��	�g
-��N�JQ�н�W�Z�[9��ƔH�h����7��<ԙ���i�XA�F_�%�Cg>ӗ���o�HO����\Ǳ$��K�l ��G'�0�����������k�(�a)�p�ǹ��<	�W^���);)E�̨j��`xy�H�m�>϶����Ϧ��f�+�2�ŘC�԰���Y�]�#	5�a����m�'�����-�"�a���1j�0ԋ�1j�Uۑ�=�MQ�Ğ����x7|���72�X����`2b�
@�t?տ��\Y�^�v�j����Uޯ�;�7zq���v;ɼ@��H�A������`GL�;�"eѩ��|2�{<���Zatu@|�wɎ��7TL�*�i��Iӧ���#�i*z�8�,>x>��s\H�y���@02A�_C��RF��Lѕ�d4W��x*�����`xJ0��:���z�f���ͣ>H{Vg��ψ�\¦�j���^���R��TU6̓]��O��惘��|�d�յ#{�q٤��V)-���*S����/_d +�!@,���PFʛg��r�D@S�d���K�l$4�c�.�����27+9�[ʧ��v�e�q���Î~�1�UP%'9sjDA��.�r��XU�4)w��D��	����V�:@�Dsx�Rz�}B�^�.S�� � RTw��qӨp<�1����_����2O+p�Ӵ�l��2�?o��Yt	��S_��r�c �v�u��Z�A-�IO��7�ݹ�|o�o�S����,���T��fϫ;� �[˧RHspބ��J"[W�:Qlk1X
�!�����3v��.B�;xJvY�F3;7�������:���=� D�d��2)]���W��<�:x�<��\����ח�.,7��}��d�}qx��.���V���0�'�;�r`���adh�z_�$%I�����}c�0:��@�.�l.��b|�$�)-�L��w����=��n4h����U��w��4|^���t��D�z��\���f"M`�z��5��Iv�y:c�~�\x.w�ۂU���)��@og�IQ�Vl��\\)Y���K[�bv��O+2�Ӧ�`죕��6A�m$^����)B)ٚ�GzK)CI�6���(�	`zk�{J�w���V8`SF.L�X��r�'֎U��-��(���r���O�:X�z�����r
��;��!6�`K@Hks���!n�|Qe[,Pb��90��܈�7���Z�D���+4 c����0�il���������8gW�����ӻ"<�i�.�YO��Q�� �+��������P��§����ZY��;?b�:�΅!���U2ˇ����6���_)X�ɩ��2��x,ќ�9�W�� (�6�mݠ��1�� �c���R�H!�0̤�G���rFf1����3�Iy��tu %��Lۮ��~�y�E��W��k{����_�b~7;��C��{Vh�����׌Y�]��J��楄��~���cٍ�v��;��}��D�j7sq�¨+�M��taP��C��}�&�������p�źU&4SOн��m�&�&)��� m)�������h��~��������)="����Ѻ��:X���q~M-���ݰ�~��f����>&wU������]1��s#����+Yw��� ��Z��尤q�{2��;Hfa��}�f�#����O(O��$
f�׊ez�5�Y��~��
5���@z`P.���+�@�dx�9�;.`��Zj�.�&B�2��CV�>4�a��VP�)�]*���X�1�\M.�G���`�n	�����:X�u��]�(!��|��^�m2;��Ӡ�3|��p/�pﬣ���������j�Ӓ�O�
�]�?CL�<?0MA�>Xd9jk"
i3�%�����Z������@�ֆ<Yw�ge���ϯNi�b�3��_���]�.B�N5�Sի���u���钰R���@{3#�z����rn/u@56ع���dG8��ZH5tU��5��?-8X�����w}���*�C����U�Q�kd�W�>�a�kU��``���=2�S|(A�~�-�-�c�� 3��������_2�����~ '-�4�9�+ˠT�ǭ$���Y��T��8�li��7`hě�_�5�_�(����h%��KL,����).6���5 �+0P@�<�6�X�X�e�+D�8�=mB;d�a̤cGn�)�n�V�;�d��c�+�Lc�J��;�#�s�û�g:S�<`��T�"�����c�b�A*R�_�;D79��f��C[�+jP��m'&V�0~I
&�3v2ku,BOO� nqu�]�z�2�w���8���(1Ì�yކ���ɳu����%��{���dq�";�o3~�Z���k���<�@tG\��xu+�6�T·���%�(���ڐ�o��(�K��x�y���`P�<�]���V��|lH)� �����%���[pH 4T��ܚ�����Du�w�0'o�%�А�M�� �%8�n�U�� C�Yf�b�a��bE;��-O\�H�-�BZ���t|P��
���l*�B��K��u3"�������J{�X���Gp���$.y��@o亏j��]��k*(��mb��mea�]tV����%�g�wK����U�^Ub�L%B	(���:��.>��雠X�� y�ޚiWEP�xtoq*#�Bb�-dOPEք��ew�v 'Q&c���/�tqX50���G?7�~j��eR�]ߺ�%�����7>Z�)�'�� ��ʝ���rG���˥Q �oZC��c���_����XG����j*�A��x�������0�;Ty������6%�jĄઁA��J�
P��e[zOZ�	�|��Ơ�@������W-�+��O7ʩ�����:0&�� �'T�p�F�:��8S*�˟*P�=o9��E����<��ق����L .ا_��/��rzj�.����c:���oes��:R�5 9M���[v�nߐ��Y�jHMm3hl
7)��Ui~����1�:���ʸ隡���H�VG����DP�x;GM3�sG�Gk��z�q�Nӷ��ŗP�p���2@]ńy`���u뗘*��5�N�L�N��� V�d��nSd���<�m<�
�9;@��'"J�Fݫk�ᣈB�?���-k��$n�j���l�ְ�v4��ԐFr�}�h�����"XL����t>���Ȍ��R�'K
w���~�^H�h���A���-�Q_k��̮�M�E*1�yh���3J��Q� &{��|dS�G_z�m�N�����^ňf�1H���,����1�K�_Vh�^[\C�#au�M�K�J��I>���B3�m����-��&��xII,n���j���Yhȡ��bIҘp2�x�P��9��_�Xb5�"��탶C9����tΰ����G���;g��X�lS4�iO�:�[Nc�G�Ϡ��X�Xi�k|��H�q/:,3Q�6K4�K�@b&�qK�)����mC�[}�_f�RK� ��kjd�?��EtN�GF� 8�Uõ݌	�<��1b�O�x�a���AV�}gi!���-I�!'OfQ�?�u���&\��z�l��bl~
?� "_b_N�q��z��S����2�-�qٻp �#��1׽�0�@3�S~�H�;�a�ٝiM��!�!�l/)�&��,	�N挜�S/��C�����eK8�����Ž��!YoR؍EA���`�����;���Ϸ�a�~���ʃ�%�5]���[�+�s(̹���J�!Ϛ��jL�^��E�Ё&���w�>_�����-���W��e�ua�c���b��$T�X�`�s o$S	^����N��go�sk.	6�hΪN$�$�4΄�N� �e��������F��C���F:��@�K �%�Q�CI�h=�x˓D����'~$˼�>������a?>�r�Z��%	���f���KTLA���墧�[�Qc���3�M����;"ֆ��h� �T�)@�\�G��Ƕ�m?�ʂ���nÕ��?�QJQg(���\���\݇��w
?���ރ��[��_C|�c�*Yȳq��`���I�y����WA*����>q�Z<�C6eoɺ��:�W{�e�j�yẔ�D�uJ�~�G��9�+p� - �&�3��P~}��"���b�V��t�����H����\S!J�a��[�Sa��N�M:K�@�S��	*���Bh�6b{&u��L�/�������K��@0�~�!��앝����}�=���p?��g��t$�$k.�����j������h+Bݠ]�������-X��"^�=d�0bO�@�Uz�󱌿�����X�H{�� �}�q�1L��6m�r���K��v]ݪ����И��׺
���a�������{��68miy���B�<��b�	�w9�XO�M��d��PKv�M^avF=��@��B4y�	0��=�\�΢�N��l+�9)��.�[� �b��j6�$�<���{v� ق�2Q#]�y�
��ŵj���`8������m�3�ֈ��V�\`��|��ځ+�w0���2�o�z�� �J9�?�7�3,պ�ɝ�CC��vX��+ ����,@ҁ�I��J}jCl�Le |`�J4�h��csZ5��Ο�
��(���*�[��z9/�����~o�}��;�|.���Wű~Yx�3msߟ�\ C�KA��|<�����Z7���A�3An���<e>��zk��W�� d4!�%�쀅�k;�����<����Z���
����񧮸M�H8�3@JIJ�Y��o}g7ym������?1QX����')p��7P�ʵ�M/,�Br(R�ɪi5��a���5Pm��e��� gKi�d_��TBIв3fcv\m�ݜD��=+W��о-�U�Ż!�+� H*�nI��D� �}Fғ�wN�e���@�&Q���ع�/Բ�E]~j�@���}8 �~�e�U��?1�&�+�4�4����͚�vb@��ֽI���#>G4`/ˈ��-ϋ� ]���c���r���$XvwT;~Wb�8;-snv��6��w)�����;�KΗW$a=l�~�E��5�`������C�����r�8|9;"���Q�T�C%A屿��?�n]�{��q5N_��-^z���o^�����%��������f��PÊ����ӏW��J���qp<>(H�(�'l5OF��e���,v�������a�Q� !W� 
U�]�U�[=�����5��JXD��͊�v�W:B�yh��c\�}#���'ŵ�D� }�~�Cb���ǽ�7J[�㿖����]��)(���`��"�ciS��w�{�!72H"j#p'�����h.3��
ɒ�+
[��������iQh=��*t�3<� @��}^�z@73+�4�Ii4E�u��eN $�=�M���{���! �\�t�T!?��ni�rb��x�;���6�.�Q�I��Z �<
�yV�z�[g���ҏ�Q�H����[N�kC�B9����ئV��ϫذ��@$36���j+��=Su�8䧠T���I����D�����K^�ـ���C@�1  ?M��O�T�%͉�Ǘ,i��鋡�!�mk� �"��N���,�2?�;8`@/�X��w����%0�7� ��aO�W����*\����@����׉��5�r�c;�nt�]��x�	�� �A�/�M�J�[|z?��������Ը�CU?��t�Gw��r�Ƙ���w��4��Y���W�l�a�ќ�&ON��'3d2Y�4��ж��sU�Z���ʖ �eO�����M��T��fw�&��B��\�rNOCJ�fvY��㖟^e�&��*�j�4^}% ��	�Op>�t���][���H�����TW أ��ZZȩo��z��x?&1S|VT������v�����w1�{'��i��T�wJ#{L���\���!F�G����ł���>�1�M���%B� �E��Sd��,vèi�'�r-sr�P���~~_"l��I�ޯ��JU����YiB��-:�6��M)�g�9E��"�>�4��t��kU&�Km�;c8IZU�Dof	�n���i��C�o;�8��l	���k+�8��i�X3��`0��`�~�yA��I�R����(~�F�]�ۡ�=9��6 Ȍｼ���'� l���F0����W�j�HS����㰩�E�> ���`N!��8pq]}~up|_$X��|O|��r�i ����^��|F�"�G�i@Mii�G�줦���K�Q�_WCd���X��ok�)���	j�MgO�@'~�[@�ʠ�0�J�C��7�"
i�ɰ]��!�rB/��#�]�Zڰ%��j�\�j�'��6�7Q�ժ'j����K�U��c�F/f��_nQ��ć���3ġF�*.�N��rL-y~��QHW˅sZ\��s~c�����=��$@GK-�Du�-�f�UX"0;nZ�:�=uR=�#L��x5U�*���%���'��6MA�J���7"Xg9��O�r��)���P�|�!t-�{�bk1��>̞��N��Y%W������Q��#�E�����k��7��_Xm��ə�w�j�v��Y~J|<�Zp�%�}��<y���A�>k��!�
NF,�#�~C��˾��ma�6�M��� ����-gy�m��\�+���~軎^�'�c\�)(%Q6��0+��L3�b0��w���3� @:N�F����DҢ�|��f��X�NʭZ�	c�E�x��ZAї��>�3Ϭ���$w�����[��6u�O0��l���	#�2"�T<���'�3A��+�z�Xƾ�tk�U�Bjfv�I��^�Y�(�*�T~�.TQ��o=!������!O\%Vvb3���R-˺Fl��69V��N���N�Z���Y�����'ǆk�0�4�*\����i�={��_�,w7��n�cCq�C�����z�bQ�sK!���i�Z~%%Oj���yܠD�^j�2k�Y0T ��O����X)�_M��Qx�.:�`��0g�k��K�`c~��.�N��%�h?�;�{�wb�a��x�,��&�+Ϥ|z�+�R�*�2���|���w�5_�N��T`3~9ԸX�V9�����>��YM���K@As���~&�1	�O�(>?@�]�z_��1�J,�ŀ ��-�|�����n6�*8�(�CO�j��5DK|ҫǮUb��WqV�͛hͿ�҄��/-��x#Y���b\�4ܷoL�fp�4�4���e�+z�cz�����a<I����Y�Y������n�
+�'��R/���GN���9%�m2^PnHU�Ͳ�H��I�E�	��m���=��b�#�N���]�� A�A��[L)���'8��� L�=�5�Μ�O�� ��'u\~y�պ.��Y;C����+l!Mn�>)Kg�;
"^�Ԝ#��b���vR�׏ZI',��=zm���k�FGxE�������[��)���7���Ɔ}��aY����"�	^D7}�,t��m����jW���{B����l;����>x��
���86� ^�b�
OC���S�!,�_�9�]�L��v�ʛ���k���sk��Ê^4�'�R�L�(������+)�=Z��Ƈ��4�dq3�B{��#��x]-Q8W����!d�T
��˂[\ص�ܕ��ĺ��V��MYH��YdZ$b�3��*#\�u�BM�������\_,�8�4k��3�!RȤ�=��J�縟����Ѿl�	�~P���I�����Y���9hv�G?���3��%&�����?H��-�[$e+Ѧ�Z<�ю�����%k,�dq^g��p`<;�VȂ���X`3����5�C�ش�r����Ŭ�~	h~�������U�
�$�fC&��.��ˍ��yv�T�KTin�U�݂�X���,�A5�)��@a�.��FKU�oZ>�8��z9��ʙb�t� UO��T8v����ғh�m�o�18��@����v�$���8���$���U�}�p	?��B�\�Z;�ІT�]�k�����{�_c\��;V.L=��=|�z+3�
On}eP��ӡ"u+��?C�뾩��O���o�Z�,���IvKƹ�\�V1���ټ	ɬ��JI�fl�D��5��5�QA�ik�Fo���=�'�5�B�%�gb���b�����L���m��iC�>9�ɇj�1�E)�~�0I`Y��|ar��}�l�0�-#7�����g��=���QN3�ƺ���k2?{a�2M�<�80��!��&;����T
6W*�R��c�?fmlսe�?��M�N^y;=�W&"o�-2(���y!*�y�z�_����̡?���E�n��X����D5�>6Q��Oi`����h�1z�s/{Sz��{�{��!���R@R��U\�Td#Q;_�+��i��d�_�2�/)f�̉�ͻ���aɔ�����ȼ��*�.�b�Y�b�����蝒�W޺E��`W�5U%V�2D�6w�-d��q��SK�(��h%3����I��#�0�8P�,��ү�x�ԩ���ĭ�#�$���5��d�1��5��`b��"r曺��/([-��B1c3�U8W�{i�qZ��|b��v$_XV���Ϭ�������G�x�4��Ս�m���AE��q��qr�?�]�`T��?|ҝ�x+�JG
%&���_��9����]��J/fy|�&>�������3N�)�F `�??Dg�����tp�Q�7��6Y��z�[���xG0!��͕f�;��l�T��Ї�Y�zKFU�O���x$�.�N�}}ۛ#����`�..~#�@��²����F
%����,�zܳ�q�y�%����-
��B��.m�d��|5L^e�웸�f�z�P-�o�:�aȄq����|6��q�z��G������"�*\��BD[n��};��p����f�)�LY��ٷFr-��ncE4��n]IL�|`��.<=D*)�.�Q�	�迸�Jw�ݠ��w���R]��G&���n1$�}�h(1��M�b�a���%_ӵ��'*V'�I�?�n�<�s6e�!r�A��j�;�5�@x*^|�/0?n���@�w���'U��X�k:��̹�R��$@̦4�}�Y�ƌu���ˏ�3����A^�R߂�S�j��,b0Xʘͮ̄2�Qp߄��k�$�Ȑq�+Q���!�����"EG�=����Z�O���m��B�iRI߃�G\���LS�.�n
q�ܼ_ozM[@Y����pL8�����i���U�o����u�ō�>��
%=�i�ԫ��#�f�� �X�	���l� �dC`��;�2mzw�L7FЈC��|�26
���H=�3{ے����+$Q��!jZ�|�.s�f���+K�V�F
��/ܕv�Q� ���i���Gg��x|�̋�E�б�/L��T>Jf�� PX��c� iQK���v�U� ��_AT^�m�y7T`;1/��Rב��)�UOy�r��������+0��_�ث���H��K�`�1藰�T�ș�:a���k��.�����@{����yIz	Y����a��7&���N섊7��뿑���&����ռ��B&`lQN��v3���p�;ۭ�:���M�cw��<o[�	M�u�eG���Q��CWX�uZJm��%����dU]'O�iܱ�����N��T1N�m�3�S<պ��uK=u������qoXԦ$�_�>L�]*��8ӇߝiN�a�@��9�p�ŕז ]Ы��җx�)O�-�^�礱c���ȠW^�.��t���(�l���7�1�������9�p_�ԿV�7�ׇ �R:��{n˷�G�sgn?i���T&��(���Vꖃo��VI���m�	L�'��m��N`y�ж#�=��E�����8��,ɡ�+"P�g�7S꽊�#�k��sX�(����)��&���Qj���S:�ѵ��E�lA9�*�|�J�/`����G�m���b���:AC-e��4�-�,��iwi� K�ϒl�V�t�ݎ^�?s} d������#��
����+|�!t�-bXP�r�e�C��	�	�Út�~�8�
��Ķ�ô:߰j���숛�N��TB%
�H�#v}�z;�ʫ(Ѩ`�Y�J��|f��O�uFB�C�ZR�lN'��f�=UJr�����S\�X�~X���5��)�b�!W�]�> �Ζ��9{�����ʉ����ă�O�z��z���g�
F��ʀW���[��b^��<�w�Բ�ʖz����"�����;��K��<���)���^�NQ��ckٮ�4�9�)YJ S��}԰�F���^1;cvFb�)���I)�� �@uizJ6&9X�*SWld!�m�E���r)R)U�k[C�����W0�-	iƙ7p�zUS��HuF1��:���b��P#��'["h�wX�Z+���΀�SH�����%cC��Ū�,��
����P�	ل��8��%n�aҟXA)���ґx�d��uܮl_,l$s��7�ǎNH>L�mz�(�e{�b��)���j���y����sAU�<v���GǕ��λ�d����f�B�_�@�_݂eǈ�q^��Zpo|mr�nEK`�a�c�Z"��R������L7ܫ�1�Ū`�A�RZ��>(������ˇơ,���!�=b[!c���{T �.Ol!���5ü���@'��>�0ܬ�}b�*�[�"�%�S!V0�{M�b�V!
���G\ܾˑ���Y8�#~��؎�����Z������vcv*��� ��]��,�z3LT7��%�Rs&U6r�G-b���|T6y��a�(����Ģ|)�Ղ�HR��G=���0uq��x`4V�P�*�q�Y�`W���7h#>Iw�wI���ѝX
˖�;)y"M�B��@�l;.�τcd4�|½2i<���j��QS�G0oV}�Wc��bQ�b(8-��qg�]k.l����E �8���硶~��d����"V~���R���ش���B�XT���1���RZ�S?ɞ�2����_m��om�b%c��?�i @$�SUl��y$��A�P��&���p��ä[�~����?i}���6b�̙P@M%`J�"fSC����;�/�1��UI-��M6x=f:��r���-rn}���
���R���K$A�`�,ھm����5�HĞ�5s=mĜ�r��NVc����6;'Z���S�Bq����2��CGB��P'�& ��g/O����yTM(HO�a?�<��:� 	�S�6��U�A�z�[�P;L�Y4��������X/k�j�>���b
�=q�WF4�t3�|���)�j�!�⥂1�a+h,���1��1O!4��3	"#}�� �f%��钸P���|E6�
���x��&fĐA�i&�!N (�s�������2ءal��c��LĂ9K������<ޠ��R��*	Q���V�����2�a��}I ��V⌎]�)���NI^ǝ�i��F�Kь��\�3���E�3oW���-:/�Jy��5Z��ω�����K�N-S���V	��~�E����tI��u��� =ϩ`�y��Z��~
�D'�4A�����n]'�A)1�-��)aS���j&$^|[�0*p]�SH}p�h-���}� `����	��3,Q�r&fIy�7?7�YA;Y'���a�(3��w7P3UH��M����Uu͟���Y���g�-�&ȳ`�W���P���~���9	�;�i�-�KăEh�kZG2�䩗�V���K:��>J�Y#Ԙc!��������~uUޛe���D+��?�Ǉ�ո��Kl�r@`|h�w��G� ?=��1yՁe�]`u"� �(5�)$+}*L���#��)��� ]��4�.�,��ď�����������ⷃ�#F�535���9˔�F���u7p����w���N�'3��4u�W5?f*��Qx{n��ʧ7��H��E���q��qX��h�s]�'4u���MЬ�u��PP�qjX�5?�%��,В	����޹x5�Y_�#^��9�+�'�løLЖ��I@KQ����`�ȁU܈S�5�����Y�#<p�ؾL��kY��j��5j���e?�����m��!9�y��d��C���iB�>.فP�Y�ڊ-I��-��(o�9=�۪t�D�i�>�>uA�U�>�ǂ/Z��.��&��|�d��V��%Q�
� 	Ψ��6�n��X����wIW�����W�#u��>!o��p�ʄ^ɧ=?�	G:���g�D�(�590���X��r�t%27go��o�fQ2_s<���cC����|�Ǹ\�`��\�`F��z���{�2S�'6a�͆�怣>�8ʚhR���8�C��@�2��+�.N�Jɍ2��9��ll����ղx̿r�� %�Q���8��m�9�A:�������3�=��
�[��Ӹ9qU�
���qƩ3��,ӑdkVaB���$M�#���<�����T�<���Q�ƛ��*��;��9o�[��S���7��c��M�4F@E��9���1��tD��İ�s:��	�R޻�ZM��DQ0t�y���cQ���H�$xsT�l�!��lT�'���Y�Q�V�O�% �ϱ?oT%e�L	AF��>�hTy��dm�!��'�3LF�ޅ�o]��:��.E� �0��mh"��WZ0E�~;�=�
����NG�ػ"�uy�y�^AZ��v@��H'	�o���������q�qKlÉhF
��_$�ܧ��{�+����s2ڮSz��`s ^8���Uh���Y⯦�7_�f,��_��濽{��Hm;�A�qO������T
��p���~l���a$�o�@�+֗+�V*�R�^�FBP��U��FAT�!��X.��k����>�^�� �\O��9�� 7��r=�0���) ��!�������#����EA���y�VhG%�ȩ�
&��HMn+^[Pg����\��Kj���|�MK7�4I��4������p�ꀸ����u	�4��i��J��c2Q�xX��o"2ʃ(�ɇ��}�`��w44D�	I`O���mS����̌G6�òl���]&B��V-�]��C��<������c�UC9��p�{лOuz�.(��=V�
F�1n�˩60yn��D�dq�cۃ�\��s�DW������$��ZU�ߧ�K��'�R�ܾ�`�i���!�>OY�������چ��_�]���}G�l۷q88J��+O>�w�7sO��D�PQ���]�4�����i7z\p0Zm?�m�E��T�XH���T�:c}T�1�J�W��퍘�t>��1�T��K �ˬq֘�ka���!�i�-�_ך(�>Z|A|a�>�O�SG2�۟o6�_�A	H�;����c:U�k���d�ݍpM��D�^��q9g����R���K�:��(4�px��F �%3��1�нCk�콑�w�uoT_n�휃O�UY�{��YP�3��!���|��5\r�.q��ZN�����LT�V��4ۃR+�q�gTzV�����.�#n�>`��]�>�_���TO��
�r�3dS���^"`�Gһ�OXs/��_�3n�+H¿�!��,��.+R�#���Ŭ0�@�P��2�h�
@\X��p���{0)4R?�V*Wa-Ϟ�����y.��S�nIv�l =�'��"�Өk_B���k��-�w&j3�S�uO���J��#��s��� Ȯ��J��l��G��*���zT���t,���eh����@l����)kЬn.�d�S���0��y��[��`��V��%t1-4|m=S�����T/��n�w(jR� ����6�>�����4��q3=��C4Ogi&B�t���7�'�3�<���^OH�225����2�����ǃ����7?[¸�APת�#x=����߯�Z>�^-Az�o��箛�� 	�p׏��Tk���qr��1��{`"��C��)<��?��V��G�\�s	���	(���޻�j�b���"���!_a6%���Y���k ԙZ�R ��R�$��m�O/��t�����K�ܽ�z����qbQj��.x�c�Cz�Ey*���un�
�e��ƣ�%Y�*8x����Cv�ڳ�o��'V��~ǃ�b�|��e�&>
9�&Q��K����5�8�+m�"��z�巯�&�2��=��y�JB�5�B��$��8}���3�*m��t��&�0ꉐ��LQ/�!�ygk�/��5޷n b]����t�ͪ\�D�� ��i���X��Ɇ��x�O�n|ō�@��&$`��G&i�����<e��BY�S&�0��3�)=�m+���]h�2#�WI���pHʮj�;���L�sN�\;���U
g?��O�G���6ó�	K-,�{&!�'tu��}��ֈ
�m�̷؞����䮲��Y��f�.�:Z�VŻ!3a���__"IH��좍�D}s�eVA����NM��ۆ�?��*��w߀\ۿ����G���uyhUo�j�p׳];�8<(��7���1	띜J| �������;�88�Y��+$����h��@u�������|%"pA�<P���6
%c�.E����()�U��}R0��Ϻ����2VE��ؖK2f(Tv�su��n�L�4����:b=q�ZP�r�n���2�݂�|�B�n�k����ꆳ�_�!<f�oMr�dv�4�]m׶��(�L��7�o���v�Bh���]�˷d�g�ik[3�i�l�=ӭ������Q�o����M�Z�J|.:�z0�'|�G ���������i`Ǝ���7��I�IQ6V��,Z#�w�eDW����ъ#��;��oY���<%G��(b(����D�f'��{{=-;��=%9�TC#J�×ļ��&���[ۇŘv��&�Ӹ�r�Ԇ�QN�j�UU�5�u�1�X*wO�����M�{t�L�2;����!T��N+���\�9��X�w�7l�����ߎ��ė�Ŭ���a�^a�'C�x�\��2]�&]� ��H��m�3j�֘�1~Ԫ%�~6zC�p�~j��,9QG1r?�ݶs����T=����HG2X��b�,��R���I&V�?��Hm~&IG��Hs���T] ��onO��ňX�2�/����7��t3��_SbUX���ee�u��4�*ά�'�W^Io�~��{��kˮ[<g}�Ī�q>��'�sA��4�>����F��y@����~T�����z��e<��k~�B!�z�Xt�.
��WkTw�h�RK��j$��lJa1��SkS1�D������ތ�A��6|9�QRX��_���4��2�G����c�J��( ��WG�����/G�d"eUZ�Ѝ�~S�d�/��M-�U�RI��E)�	-�+ �G��8Ho��%k���p���{��$s4�T��W7
�Ö>J�P��W�'#�?f��N[L����G�l�
pf�bM/K�
��[e�~0a���w`��buU�+M�� 83mU��o�����K��(?<L�W^v�Nk�}p��v�Ӿ���/�e� )w6� ��,��u܃�Gb(�N�h���1�{v��8��|�[lZ:N�S�`+��@#�|�2����>�ߗm1�7� z4L'�1yk�Xֶ,��ԥm�UZ{[��Z��'e����a���=���R���&Ȩ�����GՅ,WB��]�����_���c�2�f=�ۥn�[�IW@21���םL���χ/����ܾf���R	�1Qp�ߡ�]w����/�(A8����'�.��.��D��̢�����Q"@��D(L�؜uA�<[Z�	}�eYv��'�
P˅���bG
:X����>{��"'"���dl������r��#7vRa�h���/@֬qK��a���usnO�sN��/id����'���x��/ӥe���7�����mI^���߽�@��p������قj��4Ҝ3��J�|qY �C�ΐq�ɸ��N���C+5M���3�)�uX���HI|��S5�!����z�}j��/��ȁ@�!�-ɞ�;坼8�%�9��iR'AUin���gJ�zn���-��@���JD���Ҙ^[v&��{�mo�⻘�p��{P�b%���^�
�aS�x�Ą���"�/�H�䋢��a*ϕU�qE�Q�GisK}�W$�AvIJZf4���a�s�ZT�(q�m�[\5~^�~ߖ�V��q�T^i����
�������u�k�J��9�#p	���4U��=r&��A��|�h�	�xfKW�\��M�.� %�V�nt|���r,~��M��:�W��h-�B�"���t�_�A���=8�L2�����L����yo�ʋ|��X�q��Jwp&� �����`[]��Ơ�u�K�q<��b��7Y� �e�N�2��'n��v�W�q��|kX��^�^��?eP�SW��������<��柩+���Nך)���~0A�U׷�_������*cx�K�rH.}�V�%��������#}M,__{>6E?��d�<�	��	tY]�}���qR��(�4��VdN�7�7F)��˄�͎����սq�%�TD�?-)�Y��b7E$�g͝ ��}'��713wG�d1x�<����E��LP󜶌��5���j�/	e8' !$�I�!�8�k�H邼��5�����["�p���_�Q/�bl|�C�I����WP�m1�T���R'��V�|�z�E�������wg�Z�q�q��Q�U��6Q�@�#��V�;�*�w��Z�9�5̡�+u:8��W�W%�"��ȼm� �G�͏j��L���%�}>�6�X΋[G+�C��!�6��歆֋�e�Ӆ��v:� ��@�ĳ�ᜣ�)=��)ɱ�ϩ�r�қ^�k�B�����nP���j�,���m��lq_~��FO�;8)K��W���C����]�����ܠ����{_s!K�2��_i�
Ldm�U�ʉ�r����d�ݾ1s�et�d�(�nϵ����"�[W��_G}���<_ ��
	���2RC�J]�(Hŧ�ڠ8�G�Y긼l�B����`���?��ǥ��Fěz��$4��<����Yy��Rd�>���Wx�.��﯌b�M<�$��J �/j�Ì�����[���(o�Դ�+��Q��zy��(�:�o��`(�%w]nkǟ��Xh�cr(�L uofu�J��B䮅]$d��^��(U����!tPN�������g4��@ ѹ�wTq����t���y�?+_>w�8��o�r,���LI��E���Q^Ho�s��]�(n�(���M�R��Ѻ���OԲ3������yI#�.���ϛ�Ůd@`���#ǆ���Ss"�-(�)�JWw��pZ4��_�%��,Jt�����@�ŭ;p��¤0�*i&a�1 {�fu Rr��_dIA��n؀�Ȝ%�v[1
	��^�0u�ݳ��j���G�1�+y���a-y���*�Pά�$�	�����"��Sjd;�%n�׻Kvg�o�\�_�haR��;8Eo����e����'�T7�L	�W��NvN �,�ۧ�"��}�ܽ�o��l�Bԥ�K������s���@y8��߹h�U<K�ꦃ�*�@d�r[~��9n8ejO�~PH���j��tE�m�}s~ J ɧs]�o7q��J恈 c�aؗ���9�����g5�g+͇��]���P��٭�Q�Hy�'#$c������D ���Aw� ��-��t�&0z��p��;�a���>u k!���?����1j�-��d����H� !�Q-����5�9T�G�m/Oڣ�ln��1��k�S)�"T���f����9)mc�h���6�R��_���өc�>q������e'�]�����cLW�����.ǐ ��E�MnnN�@��Ih��h�U�B���͖�K�AOgY�E�';��L�{�xY��9J�ݣ�# ^^� �����M�a�Z�gzA)�Q�aW�DI��N/݁�� �])C60#b����B_�O��ȏKŪQ���2eڬ?��S�ݻD� ��ttM)�����b�N}��~fMR#��C֚���	��&ó#r���-=l��h�҆���@�L��a-J'���&n��>��ƼC��k��P��7��������|����z����H�"bb�(�6p�ZO1\x��i�W�{I�*��!9Q��c��\v.u��]�4��q��C�ܗ�2������e��������?�"Z!Pr�/��$�4��K���hUC�^"����T=��SFVk�$ӗ���'�O��}GfF<
ꂿ>���+{rV����3���g.�.wv�d�v%���$�` ������ip��9ڵ�;��`ڥg��	�^o�Z~A��`�,�PpE%��[����<M� ��_+
n��-#Q'N��H��xji���ps-η�E(ɨ8D�ۯ���\Q�4>#d�2���cx
��h@�y�!�����1��g��
�"nP�a�͝raGj��g)���qמJ?�Sp�&��0�yx>_�-����K���p��/� �k��0�EM�ZR����9A��ߏ��,H�*�y<������#5�"�d�&�z����A�:p��2�m��`��0��3�V;Sp쾞.a�R�t�Z}�h~7I=�w��9FpM� {+�p�!��`�2�9"04����x<o�ڍ$0"=%Kv c)�!EpP�5
U��B�~�~i�R��a�c@���0���^ע�$f@eI��ѴQe�B�>�m������1��ڗ�G��`�e��v��[!St��ko��{��-�J�E�Z|�6baA垏�2� 3Kx^{רj����B�a�4�|���毖�#���)$-u>���*c
$�O�3s�[��jF�ٰ�c���o|w�밿��3��8�^�}�L��d�<}�+���c���
1��l��O�O��d����<�d�Y�p;R��{��JZ�����m̸�m7R08�����Ő���xL����R�����+��k�4��F��U��y���@�r�ڻW���`;�L��T�+ն�f��N½�k��f�"LF|�TB/o�p7��ܗ����x�:_Ĵ�s�S��!��?Վj\�A�k�桋���1v؀S>��e��K�v]j�w�0���@W��2��4�9�ӏ��9��J	�y�=�κM�������i���՜�H+#��W��\��"G�-��@�K�wX���0�+Kps���q�6���āZ:T���U��P���v�ELo�z�ؿ�X+_�����h����i ��z�J�̽2Z}����M��^�\}l�oqk��u�ɻ�}F3��i��!�<����ɦ�L�4�ވ��3�*�1K��2I��*�VɜƬ5�p����U�-w�Ռ�̋(�s��l�e�)͟�L��n&\&YT$���:�U {W�Ʀe�$��~m?����?��cW0����p8K��Q@L-�w�X�B�K.�N=��Yoj���i�oȼ&�t��J��8.􇗎�69i�O꺢�bJۜ���j��X���P�VK3ۋ��}/�t�E��0R|��H��N�؞*l>Y��<�w�0���q�|���7kX���������t�t�ZB�q�̝G�5%ӯ�gшE���r���8A����Ϯ
�I�X�f4���v}"
���_w5���lD�p'O8��Z˯!�ZJ?l��-�NU5�ڵ;�>jttp�]y6`�,��
G�$�#p��D�����Hk�r�NO�������稠7b��1�7�	�5��g&�<�8 ^Ť��s?6�"X���D}w��j�㉛_֥\3����av��i5���10܃uHq���#GT���
������7nha�����k 1��ph��/�Ծ�����q�*�G�ޕ�V��b+>P�A�X��$���2��6�FDN�\��ڴ�5�A��oy������?�o�WE����w��f�[��〝���=�,%?R�w�c>fڹ^�6�;4,��¶o���Yϼih�m�)������j���K���߹�g�;N�]
���"��=
*�2�^��8�DS1h@�-�Ш"�<Q��RFG��[{Z�$8��y^��q���cP�%w^�e���;,�#]q���4�c���Hs�
���W-�}��!yw�L��P��0�FVͬ�:o��&��e�?�}s�R�hy6�J/Շų��9Ʌ����8���;��̜�U�c�b����Ć�Xq)��Y�r��(��wcj�O��+-]��.��D�(��˼T=�7��(r���[*6n�bQ=k�y������ZY?r�L>�O��N��K6��"�����^�D�j	�����3|1$C�o|��ܨ.��^�wO�f��k�F���$�I��&W'�i����kS��M3)}�rf#�k�k"V�Ga^��n�<��J[+��D�ˈ(�.l�_�z8;4"�B�������SA'��7hHLP�|�Le]��)΄D�/"�%�V�H�~��@�FS��j?�
�el<ë��+�K�p�:֊m�Sa�~u���W����J���kb���Ǐ�hH P�����+gG	� ���j��h���Ug����ZI��U\e�F��4#V���Z��b
�U�B��֑#�� f�A��fR��{+���c�X��.�E���p�T�E��О;&8�Ex�|���ʔO�N��i�V�U`�q�]w�u>��bҾ��[�I�d{9Imv;i��Wu�p��4Pڪ|d�Y��5����9o�t�o˯"{���+��
��������CQ�I�>�P��e�OL�ǇA�&�t�8`l�3!��Qbīv��yJjX�)qE�H��"���e�g^�J�i���7��`.H�&�#��d@�!�ly��/ʗ7!\�mǄC�t�ܠ�-�����͸�q4[ �@�0���xh��&0�S+ ���F��Ɗ�� ��fz<挣�*�8�w�8R��+����fU�m#܅fA�>y8�L����wP�!���������x�0����P�S�_�=ݺ[�:*�a ���V� d4T|�pI0y����NZ������L���]����>�L�N���_N�:���~��e�k�x1�K���Bd�G�t$�S��l��L�R]N�3וauK)0�x 5_��B��� �<�j��]������D�׃%-!G���q�^�F�®�U}�ߢ��h�CJ�������XÁ��L�]�D!�&����YS���s����0Γ�ݙ���Փ�s�f��j0k1�H=}>M�U=�ư���	��r̓]Bw&�����5CrG�J����w��ȴ���/�ݞѾ�~�����o������\���;k2,�����oÙ�� �5�셙���qa}F[�D��Csv�� }��B:	N�|����\��@஍.���1z
\�i-ĩ�v�ڡ�H�-jk���[*��-W�dw��bI��C�8�1e�K���ϓ�P �p�NH���[=��I�:p�X��=��B�qĴ��YI��[஠��r�8��մ:�@����
ƻzL�q˃c�����ޱ�:y��y���=�\�#g-��ĵ,���ڵMi�G3�}��=7O_�s0HK��qHU!�:��a,��v��H�蒴"���fx��/�*但2��g(c�N�Q^aȞ,>׿4e�+Z�[M��܅��
7MYƘpA�a來��mov���֢C('����٥�`�~�2<�_�:����듀/̗�Nz7wR
�e�*���B�FZ1i1�aL�YP[����;��hә8���H��ӊ��{�Ĵn����oe[�N�Z1�M��$�
A��2�M��ϰ��{p��e=Xo�z=)�A�ZK�"�ą-���T� ;��/�N����� �n��af��N%��XH5$�Q]n�^��KՏ���C?�%�2��}cq_}�?�"��z�V�����C��&��܍?/Q�C7�e}��x�ب�&b��v�9�F��*a�E�'�N�k�]�e�Rx%��б��˅^�I��́'���Ѳpψ��oi����`ǹ7�:��+Z��|/~X�]��#��,k�u'���+�:O{��@���g����g2�V(�Q��@䁄.�_RN�E���'��e(&=v���L�BB�:����n?S�L��~%0F���s�pb��Vv=��#\���{�l9�;&����#1 �����8%6���cg�?֮c83�g2y���[�ˠ=�~D8�N���>x�/óz1{��H���m/��y  ��*&�Ѥ}3l��$�l����5ڡ���G���wi���1�����`��v���W����L�l��Gٍ�SO�0�v���ɟW�i1\<r�a�S���x��������`A\T��Kф�ATi�56$��5�enTpC��1j�7��#0��9�n�1�/��
�� ���]e��̹5�=��=���`t#,Ͼ�-��2wmn��4������6d!�ՏB�]UD�u�\} ?��D��,r���U�L���\���K���2���+�j��	�
�Q�����dZ+l�+��5���=x<�m�C�B�CK��ӓ��%�)�O�ƍu8v.�PT9���#J;�9����U��E`�c��B�t���k� �<�tR��yf�Z�@�&jT�|�A4,��v�����a�D5�����֞�,v4�1�T<�k:���ل�\��˝���Q��~P�0~}N�V�_}w�"�=�.����{�Yi����eF.�f��y�L�ثAIa�}���ďhĺc�'v$*Bc��0����.r;����^���A{��("V 8Ţ����tg�hțMVKv���a�ywb �x@{� �b�s�k9��b)v=�9YJ"r(ڃql�7~N��c��[68Чև�JnC`�^ ӦO�P�8�ʹ����tmf����֪l�J�q��_>��~A���8ܞ�u"q#��dj�h�l+:�ż�0ٰ����ٝ��3f)��w�Qd�-Sc��z3DL��k"����=���h��}�N��2�W���w���&��|��,�k7x4��,�nBGLRN=b�a�OV���El�W��w�:o澃�1*���&��iip�,��Ýt�8������q{����O�|� �oo��U���iO���pv�TP��ʂ���p�NW"=-N0���0w~#����1'\�q��Xz�"�������Z���Z����(Z,K�����0KТ��������)AZw�a�����$���t9����ui����Ϫz?�	����dΎ� 9�¥�ÌbȻą��I�&D"�$�����w�:-
�k��x�!�w�
 ;{I��N�8���z9OVŔ{����ψ���to�O�j��iV�����=Of��^E���^��[����gf��GJ������nTn >IlOs|����]�@��/�y5؏����'K0aUn�r1�Œ�*���I���v�wZF���To%�;�y7s�hf�)�7�
�-���n�$c���#������v��'^��S
�}�i�Ap�Q	K3sx�C�͸��l�f�X!�����N뀎�j�E���H�c�8>�����������ȼ%3Ӗ�|�d9�mntw�2��N���t�o��'�\ֶ� �:��mc��r�jm<��2��T5���LD��qr�czJjo��w{�hFVg�c�wi�4Hg3�:@׹���>�`46x:��BeP���Q�t���\��m�P4m�� v%Q�ӡ����	?+�p3�*#VX��O����51��������������I�,Z
����H�H����G��`l߈hYOL]N+j�Z/�0�g$�˺z��{��Zŉ��f�O�m�W��0K��t/������Q�z��W�܅7��jÀ��}9Et�M�h����G�����a������+#:{,��Q�у�jP3�j�ԏ
o�M�����+@ Ë�E-�m������o���k)���t�DY�(��̘C�����6a�-rL)؄�z�z�-(�C��S�O�=A`�����(]价%XW�&�Dm�y=��]9�O0���8�
Z��"�O��:[�����0-�O�(6!��F�Z�{K	O#�˹����-�NgW>�~���a�S��R�7���x��N�����1��~����K�9���B����b�ڌh�G���U�ם��\�$=������&�Yq������W��
tz���d��m�-��:�X��d5Rʎ�X�e��a����zh��:R��|��6�撞����PP��Vc�j\ueash��GΊ� ?v�V)�_9м�*��|����\��9��GI����_$��E,���b�T_�ό�x%�Ȱ�;�)� �og߉eA���퓰�&l�S��cƺ�4U�}�w³[�j�b��4~�ud��cg1ݦ-�cQ�C�t��Z{v*���Ƴ	�ZҠ/�}竅�ꡍ�h��s�"���I�@/ޡ��~��'<�`bD^NR;�B���X{vS$Lh�K��d����k�����/o��Q��%?���0��I5�16��؈8��I80ꌽ9�ӯR;�IA�OM$�%���e�rS��H�s�e�����ߞ�h^/�Alɉ��3�Y�۪����A�z͠˵a��YP������0G�<�J0�mݫ܏K�����@�����SrFQ���<:�y���K�5U}��5��y���%Sxh�U ���ե���1�s�7R�v�*���I�V��%�*�o4�s�!m���Z�Tb�Qdk��!���3a���B>�SD1ך0��_��3<�����A��5�N�=&�$mv遰Lm@����W�C��db���RDy�j�TQG}ݵ���6�wV��8k���E�Hq����_��Y9߫�_�K��s���7��8#d=�����.�{4�U���eϥb>�����������>'٨��O�4 �I�bB������c��>�B���'�����ي�>�o'u�����G'��[B�e�1�ޓ#Q��_�|��m�ꤳ�v7$A�7��{�]�lխ�~�DAُ�&���XM�A~7�u�u��>5+��%��-Ǻ�S�|�Q��	�������LN�~��'!�˛\�a%��4N�F�H���M9�At��#D����Pf>hti6z�r��\�@�sA��|��R^��Wj�/p.��q�!��X��̏�h��b@�;�P� �p3�M�D��@P�8*�����:Uʊڙ��@�M�`{��0�D��w܍-���|��#�D]d���ma�ia��`�{� Rg�05^M���L�D���^�G�4�XV���oa@�[�I�p�|��RN���,�{I�O�5vY#D��?���B�k@�.�2<g�<SA���Bm�SS]�B_v���6���b�=Rv��o0X��2˼���'eE������8f�w�ٿ�q)0r4����Ϸ]�V?k���qȳZV� s��2f�N���n�@}�ɟ��-�����Tm��1(��9ȯ�,�^�	g�څu�3ҒHVS�w�,
�t�����n����N;�����O�R�4��;�\���g�v���#�	��/9Mi��%PΊ{�tO{�f��@��-Y�,,.8�Z�A�$���e"�ʸ�TJъ�m' ��Wm'zm`
0 �(f�d�jL���1���#2�zȮ>���H��DLw���N�tf&囇܄�kV���R\�����������	�7�O�/l�d��`#WV�����/�!׽bi[��ʟ@T����a�ʢ%�y%h@r�pg�<��{���J	�[w�٣�x�����+��x=!���NE�2;�4;�;��i$m^�֖�Iՙ�4�����Cș��D�� ���z�����zt�h޵�P;t{g���5�D�	T��po0yB��GD���$�p�M����M�b�����^����`W�x5�W����'Zxq��g�z��̩� ذ�ޘ�ۇ��4�����MW��YnpK��Yv�o���n������sC���VBe�!P�K����x|�h0��A���i.�^U[��&�a�_��W��9b�V}�["�Τ̰�7������s��E!�ݙ9 �9���1�o��G�p�_KU�a�߆9"I�q��n������ԝ���	,P���w���wc�0x�%|zI�(/��J*f)�����k�#̨���IXT]O���$��<݇QU�Jh���~��a�ϸ?u���+�ʅC7q��E��G�z�!j�l�d�������"���s[���yOM!#�ʴp�F!�xb��k��xǌxJ K͍�R��\�����,����do�
��ѦCIQ���F�=����JG���λ�;Wk�H�x)�s�X��o��L�ۨ?��!ЛRPK?���{;YK�G9�'f�Q3	��V���I�r�V��˻���CX��0^�!�(?�t-~���ht`]�<��D;���ih�6yP���{+��P���H{���ʃ���A^yM�C���%|��8"E���(P�I^��*QJ@��Ց���ഃp�9�T������g�Sk�������܂�{#�+F6��d��ӛ8z��b3����2*���O���J ���@�U[=Ss�x��IO�͕�DP��\l�Cx�_�dQ�T�74`g���l�A��C�&
�����W5���>�)y��n�<���?��*�S�ӌgS\i5�\֖ZD�l	��:B���%4��]fF��U^ӑ@�H2@B��D	���|}�$�N�⬙0�"Gi�N�y
�7�i�[� �r��k���5q��e����e��a=��<�Z
�h#�[L�7��f��c-벽L�>���A��&�`R�>�!��6�&=�F8@���
���=����E�u��b�����h�b����㭟	~�hޡ���0���P���h��hڝ1Fz���eA��7H�����I��� ��R�ѸH�=����t��C��6�}��y$���5�O�% C$b��9����6�cS�I^�Ț�r:,�x���R�W��
�-p�����%^����?����M��������5lJ̵Y����}IfX���`*avذ�t/�6dˌ������p��Q� R�6�n�%�����o��@�FOy?1>s��'SB�L��*Ap����l�`V;��-�B(G���t)��q��N����ڤy!�)�i;"ydE3bb@�R��O� ^������PkGR�����˼���dy�R\=�7s�W)�!���a@��(��8���M��_m�:�Mc�Nȭ� q�u;����kS6��b+I�wX}���a����hhv���|\���bd����T�y���h����t�P��cv�~�(IN4��~�+������5	�[��*p��\���1(a�v�=�\AE8�ￇNu�����*um�5ߡ�ᅨ�h(�/٭h/�9F��*����cBT-���<	;����"���<S[ޝ���V�bt���xP]�'��4h5Hmq;y�E���
,'z0�%���U�~e6�==��}��t��P�s�;�W��i��UWO��M���ٶ�t��A�1�����M~�b�>�8���n#{��xI?򞝤�E�JF(J�6�Ƴڞy̽�(�?\�����[��u��v#�C*��p�)��yUT�-r�h�,�o�����,�|�^.+sG��,+��7>w�ru�vb(�F!�(���{��ε��b�>5��6-�TS�/y�	��i����[$�4��9�M8gj~~ꋐC�-
e6��z@gy7'��d����
Qu��-�£�C��^�$N �\)�O��R�9D��yU���a�������VY$�u7㽘9��}�;�)����hX/|������
p52�9�G�k�;�x��&H證z����fGd?C�V�Pz6��
��X 5e�i�S����/��ؐ�\�\�$��>�<n^���J��ŕ�<\�qnu��M��x�;=HVWI�&�Ij�Me�,���N�����pL���I�~`Y�D�v���k�_AE�%q�W��[ԜN?�4��o��'x�9�/�������a ��^W���U�=��n��1�&MzY�ϡ�"<Ic�8>��p
�Yt�'�(S ��75U�(�!ͤ�l�.���ׂrYYi��?��P���'|@�6�ȟ���1��H�Eo��KwS��Fh�7��L�3;���ȇ�à��e�5b��3a��QAjឤ?��a���^��N�%+����^�+m�r���h���䓬���tNfv�wuw0	�>(���"��f��%֗ꝅZ#�ƈ��	���<��1T�:+l����o��P;kEڬ,����D�d2���)�=�W`��H���$,���e(��BZ�;�c4 ��3��xlڙ.�=1��~$D�bOi�d�p��0*�ь����r/ِyX\eR���n,Z��1�:Už��No(a\��K�Juo������Ve*��3��#o��aٚC��F��H*p��Jk]��ק��^�X?c [g@a��(�Y�����qg�i�u0f�OYYi���ug��1�w8|yH=dt���U�����q7<�LC^�GG_�6�[��{݃m�����s��9�3��1����h��ZS���2h��Xy�@��r���:{�N����`���=�>~���i�4�8�wR�� @�f�_�mIu֠E��2T�̏tRF�L�C,Re㲯E�8h���}� ,�gd�J�c���f�{Q���PP��/J�0f��ůS������k�:�v�|2�%����ʨ(�,A�#��V�L]^�9�!��j`/G v ��^yU9�g]��N6���5�,�7��P���Ɓ�4z����ߠ7����J�=h��|7Y��q�m�`Z�7e��5�m�^%���ݳ�}?[㳩��V�O9%�d�����j�h��:��-��cSB)]���9^x���oBn����O+n��E�}z���1��M!<�G`!��V��2i2�πA"���q�##�Oz�S�en��J�� A��ġ�Qik]^��3��Q�����I�G�HTz��Ʒ�X����l~�WOx�
�N�f)�!O�r���^>���1��B �F{�6�	\$o���vL���ղj������&�iX[)sv��ƊF��[7G�������\��T
��j(|�����p:I��A�-�S����
�f�	.Rļі_���U��	J%X^A�F:�&��2�3�&Q��[%�U��=��E1�f��m���+a<�WV� 5�����|�L4HϏc���Y�E�}r��o4z`��D�Zg"pɷ�?x&��m�"����6ĺ���"�W�ӈ�=E���@o��L���L-V�pj脮�bT��`�5�vV�D��t�[Ը�X|����!�/}�qb�/��ES����o
1������z�+c+!J:�ߔ�_�OHv�6��q�*�����*a 5�ƄIhYqݑ�3�6�5��2hVm1��K�4�
���\�JQ���y�H��-��\wj~ዺ� �s��Eteϸi
k��i�Hc Wh��)	�w��aǘ�Ƿ��+Q��(i�K:�R�����a��=����CM���\���W��0\���D��g8锣_~�(��$|M�~�Oo{�z�vZu8���Bm0o�-M$�q��XDM�mm�Q�=k�`��QP]�(���no���)_��%�}2�,)���l��08��_�j���ڃ���9��[��ՙ�*���s����-��R�>hA���k��c0�<�M�4��{�>��Fy�V��3���ՄHX��C��H��|���=ܱe6�ڍR2o��A=J�t!�䗟�A	�ʦ��9�!�������n��̭�`'�ux׺�0P(�+�&�n7��ջ��e�(��T�=��a���V%e�Y�4#j����[���&��,�\̗�^����xo������C�z�t��oq1A@K]u�����a�rE��WUx�v�^R�+dRu&8�~��_G���HCP���ÒuiS��dIZ\1����r������)9'����  �э۶:��	�=N\?i��nI�ɝ�	�!p2�'�{m�3�Oך�D{�Ո¼�N��c���9R8%S�93��9i8;��s����t��+i>���h'Ӑi�Z��&���M��OLX�Tg�d�h=U	-�1��
߿�YzXD"���!9�Lھ����`�q�n��e���kMR9z��L�����1k�5��p�E�h�8pi��a5m�w��i]R�[c�I+��D��h�ĩ__�1��G�6Pa����L$�����������i/Iݕ�V�2-�3�)�7ܙ�y���<�Qw�a,g�xI�["��&3F�$
���A�*Q;]�����yUS��r��)�&�r�`@>:q��9���X�P������3�ԟ:��_����m9-�#�E���c_qHn^֒��8��͚e	H�����%)�ª���K��6l��	A������Q�����j���A� ~��_�<1����6ڹh�J��K{��:����y��xoz�]=a]"���L 4��C�'btZA7\t^Y����S��e|V#�#����T��l����	�����+��>���IZ���v���c��`�h�z��ݥL� J�/Hb�"{���co�޻.q�n�pT\�9DV�#�'A�il����(��_�rZq���~E�ӆ��߇<@p�U��&%a� ���_��/�9%�|<�1�G��6P�u�cp�����z�����Ef��[�w�M�gʓ�=\ KT�D���Jq�<�2��v�d)زzT�]:z?2�߮�y#j�V5|�ԣ�@S=VP��JLJ��9��!r�irD�m�3lfc�W]�����4+߁�/�eI*��N�dC�Pe㴧�U���/{�P]?r�|��}b�v&&O/�|�H�s��/��H#@XW'���<c�"�
{��9X��,�K�I@	P\�!���sY �_����ԋ]"� -�E������jG���d�! ��+Wi��skt#H�qyjO&��4��-����L���*��$e�5��}$a°C�Qg��Z��Z6��A���n��<���쐳�h�T@��񳴢.�/��FP)�קA�v�����W�H�G]�)�J��l���� �)�b��E܄{y�8�5]9���	�gm�"�	�q�[�h�O���k�<��(���bs�뇈�{0�E��c�Dfұ��܌�CaV>��
������6���>2��

� �4�T� N7���;[���S�EN[�Sy�
�����n��<��������]��ގ���u1|����m����B����T*�A�P��mr�&'�敿�<�=(��J������lH�5��T�_�1n���F�T賷�u��Z���y�'J��ȘQ�"��8�ݿ�Un.=�����3�m���U;���3ڴ�e��YJX�����(��@��ZZT�Y]N돡�����H=�wn�\a���V��� ���f�_�>uX:���a`�Y���_uQ�����P5�%��=|���������t�y�Z^>����~����^�|t�f)(�a���o��X�˃��n���H�� �Uɪٯ�N��t��B~"�_���v�:���b���Q�5�;-U����}1qL��L�Fƶ��'�39�9�u#��,K;���`o=�����Q�����`'8���A�`!u<��b%�,�^N�J�I�k�2WЩ���bpw#�x�V���� ���%h�z��+CD����Me�������Z�����`Λ�4ݸ���l}�R�������y�>�6���I�����6X���6�A�r��u����>�[���*�@y�nai�z���E��1���N�K��~~�p.��u���H�CR�؀�G���8��p�Sg��+_�b��&L谓@ !�O�^\Mn��Tӝ3�dI��΍!�t�����b�1
'��6G�?�@y����k��|�-�(=Ɵ�{z!�5�=��\�^��BQ�]cP`b����dpRo-}�,Jo�eN�6��*�0���~%@�
��|�=za����l���������"Uu�J@����I꺧Ԩ	W������ӟ��(�l,ؓR�cGw�EH�ۯ��W��f��[��U��������o���Jup��ĈA��q�M_����K�dP���>�ҋ��:i��㣈�������i��:��V��x]���0τ �o���h��X�om=�Ǔ��(���_w��p,bQ��[hS�b�_J�/�j��s>�hÅ�CITv��(-si-�f�Jk�9]�^S7r�.���(������EՈJSU��و�˩�&ɂ�7�}|b�}R������Y��sK���HC�PpxbXf���
:�$�Qq�H39���9Y�I��MNP2�Ii'�X��̈ҹ,eգ����;XkY��[jZ��{��	S���7�6!	�����6�s�F�������/��� )T�X�����'lmO��(b����A \�Z`d�d�1W.�םm�������%C�q��3�U����c�;<l� }x�	^�(���:e�"u�+TXw�Q����eQ����-��#q�Uy��H�r�� �H+�X�6��cS�4���
cʹ,��q��,u<�%=��>	*�$<�_���������v���F�F{=�{�#��,I"� �ojI��zh��u�X����'6����.��f9�L�,pg�����t����=���1�r�<j���m�AX,�	�P�����o�6 ���框��wm-?�3H���.Nq�G��K�;c,a����--IG\�c� ��yh���'�o�fMFb�}��Q��n�{��8ְ�2�'��-N��Z4Q�e���t́N�B)s�d����3)���_9T&h=ƶ�1��Ԣl�!��l=]\k�|����S�H2?|}ށC�0�\)�&ƺ��H1�&N���9ih� ��<{�p�1?fֹ4ͥ��X��y��ߒ�ٜy}@g_jy�b�Qo8���t��1����o�4 (��z���E�W�NΟ~�U��4œ��M|�~D6�c�;�l��FN�5�yB�[��O�o��\��)5��,q۾�� W^ɷ�`6�2�3O�&���	�Rw���Ф� ��_�-J�6�~E�,h��⽎�T6M�_a��\s��"B�ڸ.����bUTP� ��w[=�:8 IB�Vt6������ 5"$#-L%l�g�@\]ݽDX�o�1lL��jA�6#�+�a�չj��M�������s0�ߢ�4xW0v#c�i�Ҍ����[���l�9���8�|u���]G����0���4	�>���Լ�38)�VX�Lq����d0A\px�D��t b&�����
�Z,Ů�罈їl�{�?�PR;��:ngq4���0ow@��������Ez��Ȟ|g�\$�������@D�kL�O�BX�*�^�7p�ѯ�8����]=JB�#z�Mք�=Mʢ�'#-P��8��~�GժYS�׾U�D<PJ��Xytat��c�)v���h{�5RVt�h��&N����5(��1�\k��!��+x��Jrd��˕���v�\�v�+F�
�� A$s�V�������0{���a��0��G�Vʤ;K�U��;�S��i�����0$������'U,]{c��.3���������6-k���8"��P�i��(т��g԰�ic���sh4�B)0��;c�R��]]�5�r�� �?�����[p�����&c����~_t3�T�Ot�U��BN3~=�>g��:�	�7�hQL��Q)Œ2j�B��C�I���pE�}��w���a�0͆�9<��2=;t��p�Ff�2G���4�| ����k�1�������i�
�=F��z�T���G#�����T�d��d��J��S�J\~Z�}=�Ύ���kyv�-���U���Wq�ST�$A�hp�*��8tZ#��Uֲ�%Pe2]����aird >�/<���X�J�:s��4k4��Ց��-�b3�[�l"��#& �7�����Z�eaC��DܬG��.�P��l�}���a�s��U�>�ŠEɕc���GD����t�j�z�,�@�����BBמp(!�+D���:滠���xyHDk�k�~	dI��6'p+s�� !��/Ĭ�RL�#�������T E�6�R� �R0�\���e��D�w&�M\�9vX��w���7\�w��tܬ졘��Giok68���?���˖�BF���2w`$l�X�,x�wU���xJ���따�E0�X��CpN��������a�p3����*ȩ�8����I����W!��IM��H=����qIϫ��d8��Yh��4������g���c0�#�
�t���?mRZ����9C���b�-�Dp�ꪣR+��j~��|5�T�ǄUZ����81�k�N��,��Y�c�`|�T����]��Z���7�L�R�<W���#�o���(���TI��*��e��!�<���P e�� tYp��:��� ��u�ze	Y��c0�2��� � ��ۖ��U��:ǆ֐R��T��z�;�ߖ#@�(	/���w��	7M��+u�BW:�r@��'q��˘�:�ڲ����y�r�}��Ք���̨��x'v�7'ꉰ�RI\�i[$�L�Wb�!��[�]LB��_���+z����qt�w�չ��r"(p����M}�+����g�E��<��[-EyN�Ź��%p� �[��j��R�
CsNV�� �UkAt;���oF�fLB�o-��5�õ#5�������~���ZL�W]	<+;&5G�I�跺����'^�5��h{|��'���BX�U��xr���d[;�h"�۰OV����5ܚ�¤jgoa!����6�t�u?j}��чq+�O�T�;��P8�,�
��#�[Wу> ��	t\*6��;$Q0&8λ���@j�����iD^�։F�t�����1���8�p�&i�K*k0��Yb�nǤ����O��#���3��Cr�&��U�\,��G|ƁUI�$�zn�6���G����v��}���)�{�e5C����@��˟~]9�/�66�8E9�9b�Ʒ(�_}Q�B|�;:^M���@��Y�9�hW�h���
���N1��
�5�����8�g�&�`�&�]7y�����~��:iK\��p	�mcpk~�\���uR'(iк]�Zx��S!p�Ҥ�����^�������Ӣ{<�n{F�u�g$��ڨ~YD�=���t�!U/4�12�����y�"����%�P�R)�/�b���k����!�������W���ip [.m�ԙ��8�ݪ�)_���^�?d>i�ɻOY~#-/+�Fm�7_�M���?è��g�j�|�&��ԁ�/�48df:opK$������i�S�V�c��\T�iF�#;��+���i�6����7����w^������@�6�.��̯��Q�QR�+��k����.�ڠYޜ�2��*{��p=��I�66Fm�\�d1!�w+�u���\Ū��.���z֮`C�N<��PYti�L��6����jT�y���ׇ��͒�v(aL0�-�p�_��{� MO� ��)5��Ty�#��ʒ�ƚ���_UR�\Ř8��S3�N��<���]��2��%bhi�ۤ��Èϧ�O���䵛y���R_=�jv}����� '��=�c|U�G˜H[�nj~���հ���0w=��Q�,ؗ:�Zo?q���3ڞ�i�p���^��5`tn�uMb`	�Y?���=�l)f�M /�FԧM�y���օ�����̺�=qp�Q�"^S���y#��N(�@��©�"8��x�B�!�z:H�_'F-S-k�q謯�A�p��FVw_��|n ����W�B�_kOz9��%d�g�W�ç�>y����y��a��&3��>Q#I_���&��;p+@�&;Ӳ5٧TEs��y��r/ԑ�H��:9��o�2�%��X7'�FkX��&����Vt�N沣�i� �MU^4r����:�<a�n��.h��JT~@3��aOCؑd����֫N�օ��v$�1^��Æ�S���:�W׉Gw�X��h?��Q��TC�ziS�����)�������Ĥ����/t���M�t�w���r�K��v�Wx�n��^כ�h�*1���W��2�_�(��::@1z �ת�3'�����k�S?���<_��Ѱ�5y�}94SeY~J)���6.����@��F��>����鲧]�U��ۣ��5���S
/�[�Z�,�|{�6�G�K1��Sq�V]z�|f3�:��m�H���zd�ԝQ��6g�_���=���;BsY�H��a:��Z����b����)�L�1G�1,��7[->��.B�^�GV�0�a/�,�R�A\�0v`$z��6���F�q���%��pufv���v��jb29l`�x�tGE����Bm5>��1�{qC�m�c�և��N1�?��6�pv�Æ����-۷?@�Ӣ�`\7.m<��	��E桔�F�
���}r�*�����%���D�6����4�",B���L��-��=8WX�n���){�j���,5��E�m����е>�2+5�B���� �j����J��8t����%"�1_��%t�Jd�i!,���$9����فb'�i�+�3�I�uގ�$��$�
��l^�A����U�_G������s����:�m
�#�0>�~��T�GH][�x�i1R�l9��זC���b�NqiRN��eCN���$�<¯��K�:>^+?l�2�HER��Q��2[
h�с����^;SŮ���/�[f�����v?-�'m�ߘ�3i8'�-�1���U�oum-@�wy���
x��>�Z����<�O�}=QN�|~55����QR__��Y�(�J�́OT�c�\�U�)�h���h��Y
h���)G�+�!"�Kb J�p�\
Ԍ���S3"�O�B��G�wa_<��i�:0�$���Ź(�D��Ƽ'��uGquC��Рʕ0�����m�+1��N��f������t�TY} �#c��{��mg�椰ya����([wq�w>��8�c�`LY�KK
6>�� �̨Zb��Нk�M��h�z6�<���j���R"u�V*�׶����
Qsx ��^�P�@��1�W$�S�s�l���&�3ѿ9�c��M��5��Y:�x�1�N&�7�'�?���8$�D����p�(o�4F��d��W	�	T�]�xg��<Z�gaF�K�u �|(aDE�8ԙ/R��܇��84��FMl�� �f.���)�0֣׺�Z�(��A=4Y	A�&����!�������S����t��2Z�鍱0UoqM�U&��:2;oY�ES������Q�����(�e�;�<��B�Ӽ���X
���96�M r�~r�yK�c�hz*�s�Бe���p�yE��Vz�C��5:�д�Q��ڶw�Q��qߪ�r��i*��T�����%d���J����M` K|�opv�=�k��8�?�X�b��X\�L(=4I>4�R��!/�BXZ¯�$�{'z���/��I#��i�@|��H�1�@䙗�OZ�O�h�������S��C���={"RC�_��UU5^�������3�m��J���xc��K��"�oJ	IY���,�� 9+��� X�+
�5����?�~S��Գ��i�%��#؊O뾤�6�އ%�H���;9��c���� ����%l�ӂ�R���e��^��i}��*{�4���]�z�{<����]�0�?U�(KM<h�Q��
7aw1�rl(�f�t��#��b���t7�f���\��{�	�怬��i@ond�c�����L��W�����M|J9!,OHgX
_�p���7�e�6�"^g%�EDq�-�f���&�h�����8RI3(Q�Zi�v�4��~� �b~�`�X�ޏwHE��?8!�n>U�Nq0-@��>��Y��<��]g-�9�eW�є�z>oe��+z������$y�b��\ �S%*`�S��ͺr�O�l���+ԏ������
+���'���K����<jخ$����}9���������rY��?ſ��S�e�M�v�e^����ay�lB5[��;���B7�Y��)0N�y_z2S��1��c�؟З��c�V$ɕ\�?��'����j?y��P#�J�
�]�TqfO�=�G�0�)�Oa_�m��罦 ��5y_s�{i ���o���F<LK�8+3'���T���_�p^wӢӬw;�2�Kt����X��F�>+y%�WQeVKKA�>�%�6C�"�m%�s|�g�z��¯��(=ݼ[�1tuL�JV�z{�'�&s���o(kTW ~���j36I �=N&3)����)�� �S�v{�P]�kM
r7#��C�xj���k�.����<��x.w��e�e��)��}L���4�x���.����b�~��%�f-E�89�=q��	C��y��O?� ��� ��q_ӄ]ˉ>ҕӖD�҅��#:�?S�Q#�$���yzhD��uhSbJ���H�$��򄖖��̬.�E\�Fk�~A]�U,+�A������Ö�sL����?�*<f{�{;�@��g�{��pK�+�5�b��\(i�%�y�2��@:��Y��Z� �L�["�<,}B�=11����?������X`�ީ+0�]p*w!�vLřW/'��&R�Q�vX�W�5��1{�GQ�%�c~��O����Yi����C���[/)f+���U�t��?\`	��
l�}yJ;UJX�	��=cR��O��f4�ᠨA�7.��L
z]Mp����W����������u$hz��ɲ�-D�o�D�I_�N�����	#	T�},��}3��O�,�P�MR����%I�D��K��G.�������O�O�_v��y)����X���>�a3��e�j�nXZ)p��/��=����g��Ragv��*Ҙ�O�1W�|�	�O$����"���WУ*u�l��<$4��Wd5j����Rڛ?�S!]5w����]������#g(4����3�Yʥf�
��.3����*"���\R�r���
�0_\��k���$^��{�]W�ג�Fxb�*���@�z���N@�5��F���������p`�V�e��Є��c\l�c�%��9
�v�R�}	�Ic�W�x��(��rBD���?y�+�7�-�kr�Sb8.=wm�0���l��f9׶����1������Z�x�r����?�;T=%~DNm��`fAe��~��N�!�o��0���-b<�VE!��;F0����YWQ�0��_|���q<AY`�k���'x4�|Wa��ǭ�&{�<�gh�8j�>��+���)(�rPM�9`_�}�cע�1N-s�vw�Jn�E���<�!k���H�O������p��̙JR|���Q�j�ނ��<�6�x+�/���`�����G� ;~(��}Y��UVInh�Q�v=FN7i��M��7%$ Q���j��-fon jIpՕ�)�>���юE2�E,Y~m��Аlp��ĳ1i�qS�鴙~�m2+��'�K[�J�L�����\ql�~�1��[v��>��M4�?a�l�(W�ʲT�]iK��H�E������2Q���0λ
1J�A��4�{��[yz��BI&�@Q���	�]O�CfJ��B��mt�A1����*V�IO�I�&,j�'��֨l�6)Y(5)��>#�Kv9<LtZ+5��{��}&Kf��H��1+�� ����¼��60Q$%ʯ�\���C_49�����!���b���fN��2'�Ǽl�ޥ1����M�"��������κ��gH �?�:ݍΥ��4)�<�	��x�d;$lR�i>ƍo`R��D(��q�Р]_����GIqq��<�b`�����)��/�i�Y��e�W5fI��=��*�J�8=���FE�~�����n��<��Q��]4S)�������K̭!��W�	��ZV�h�h�4��sU{�gP��o�*��7�10��J���]t��Jb�dx��!J~��������K��>/n6��M�3���K����<�dZ]mt:E�V �V��F啰L�i����,��	E���k�GL�i�v�j���J��+��\=�����D�fAsE��f�l��8���{'�zR����i�� �1��G�u0m�I��W\��u�����ĦM7�ᤫ���/L��w��K!F�)���ɓ�y�s�����G�oR�aɔ#�C�,h"'�0�f�?�ණyx3~w�;=P2o�Ep���X�L��ZR5NXq�pHء+W�̩������{e�U����׵m
����_�7��u��zi�IQr�:����7{>�g�ң�|@j��e�_^l�4W6�Д4I=�9a�1�^��O�兗?7�.#�|�џ|���Ƶ榫�B��UI�ə�Y��}��Vk��ܲ��D����s�&�XH���Դ�%�߳�>��*	F��L�bd�i�%R�H��@�/``�Z���l�vJ*��W�6[\�F�b޴}uM�&Z[MƉY�DZ��lH{��i!�)
No�Y��C/무�UM�ݢ�<���{儁�Gy���b�Q�v�[zĤx��A�!Q�T��O�#��B1�m�XI�)��怽5��63B�FP�'��eٜ�/`�ϊo�o	��$�,��b\���30�]�e��f'7ay@�1�J����Ge
��i)���&�s�ȋ%��R�kƷ���%^	-n�*�����	P�XŚ�Y�]�NU>Lc�\]^�W��Ń�	�C*hnS���FS�D�ܪN����r���lP��),H��7T�8Y�{�o�L�d�W�����LiW�2qU� $����۶�b�_mC \�r&�p���X�����p�)ag�g����e��z��ܷ�ID��O\�Y��F�Q	-���=*���r���n�	�/C��/+[���w�6��M�3��	�:.h���D�Ԡ;��o�_��%�t�'G�9���	�mE�m�H>kC�N.Ȫ�|��H��e�S��2�St)sd�yާK�4>f� �-\|c�ȀݢZt��3�����7�PC{����$d6`�J�$��^�@ -���5��5�����ڭ�MPv��Q��`��uAi"�Z� ����h2��JYH���0E���b��%�{	r�u%�H����l��z���#�A�é�R_P_���$��U���^y>��%���Z�̌�=����%��Pk�H!!���S2C,�s%���0Y,"��,1C+'`zN!��{�$�56:a��W���T��SV>�Uhkyͣ�^��^��}7�n��;U�Bɛ_هQ��m � '�2���l�&��zt�V�y�pN٨���V�7�е2 �?h#z�+����wdP��=2���l��?00h	���jFP�� >���[��1gI�&�&~1t���1m5����v�PK���R���\%�@j�o{��O7�(}Lw�9J���3���X��k͡���B��r?葌.�8`��S���)f 
���U��� ����s��cO����Ơ�>�a�AF�g�"���~QU�(�Yb���BAY��\F9�a�80o��D�W�΍��C�v����.=Z��PY7��<L`�&�o�a���ZVD���:ʊ幉Z����ޓ�`�X� v	��������#�9v��M�.�r�栾�M�x�NE`��ي{�U�u��uY�=�9-2�Ϳ��@Bؾ�<�@��� �n�	&܀\nI�*�c�6�UC�����\o��
 �-|._�w,�~՘H@� �֪
�x�F��ӊw{�Ln*����¡�#/�4��ly�;�l���$F�t;E�xTWA��$���Ds����_����pc!
m�����FV#Q���R;�/�,T�*yٌ�)t�=�&w�{|���`\�!c���y��ِ��\�L�9dp
}�I��Am �e� �"��<�G$��b�w�����a�Vtp��D�!�r�:��$79u@R�`�-#I�һ_��:	1T ,s��V�tY���Kp?�~�s�{5!���Qw���zj��zH���2�<|$���	Ѓ�.��L7�]_@V�4�A��'�c��螠 ���ΐd��� �� (>�����۶#���%W�0��'���&-�lp�S�oY���YJHoׂ�)�Đ	�vqc��d���1}�HB'�{�{������+�$�
��8�w1��7��t��KLcd4�\��I@V�H}��}!"l������ �3,a�L;>0\M	&��+E"Gs��´��J]��S�W�s0�P�������9̙���;��}z�};/|@����͊�S��Syؼ��ʋ!�k���V� `+-��n��@���_��F���~4�U\9	��2 Jq����._�����p@�Yp�i��G��t�h�3c޵��"XJ>���C�tqW� ��Q� e��4��#=����a�|�cg)�ٛԜ�[�L���;'���/w�9\�l7hc��_�)\I޶$xx'�'�I:�uN<h1)*V���c`�=���zݭ�.��Жw�(q����%|�~|}�c$��o$k����ʀ�@x�_ǒ��n���9�(VޅL猣0v����l���aF���s�k�Y��紵7|��1��6�P�OꩢQ���kQq�q���ʏ�lf�r��,�|{�|�����@1��Jg�8`z��TAp��XD�A%��ꂎ�*�zp�M*�\��G�^��ЂO��*G�´-W]��{��U"E����L}���+�����@�k�����[�})7!���4�sP)Q�c��rw���g4��5� <NR1eM�؝�w�����V丛?�<l�lt��p�7�F9�\��`�ʝUt�_]��!�u`x�Y���x�p���>7{H�3��3�ڲ"S��#߼��q�f���*fhI�ҖM�� ��֤f��Z]%[������Ե7�7N��hy/Ȳ"v})�����MR[��3�Q{3ֿL�.i)�R���v&�"�ט���X�'����8�� ��T;�*�5�J'@6�WܷnO_ʫ����a"��ZߘBOrUU����錎[N�݄����A���0�p>��dS"h�7N2pss��nE�����j�u�4/ͬ����a5j�^��DE%�u[��iVi�� K�	aϖ�Vz������������I-�3�J�d��2[��]޷fa�|Jl���l�s����E��^u�2a�ܘ���;�� ���!?�Z���.�Ϻ'��=x�몊�M5�^��1�*4^��Q�l����p�Sϟ9���y�U���%I���c*�fH��H�nz�]|!j�͌�����!f�K��D}�M�7�H�5.v�A�Y�9���_��o3id�"Z6��f%HzZ���5������IU�^7'��c�}�EQ����r.��\Pq:����xp�SQq�t���@�s�#0[�u�N\��i�H����uXQ�m��!�}������:e��Y.�6�O�-Ƶt�)�k�bxbt�Iv�F��l��^Y���M����<�ׁ]�������]��^F�W���wi�[��)���,�fGd�+�E����8X݃�?��bYu���N�X��pm׼O��a�feY����їʧϳ1�lo��5f��mE"U��/��>ϯ|��W�����ı��Kh�l�d��)�5(�.����	A<��7�qy��bI�n�ʲ�B�>Y-{z�>�F����)`I���@��p߂��i�����f`z��6;v`����mg�U�������	�n�1Ν��r�o�3��R��>b��(���+wj���!�gb�ǰ�O,3x�.(=�63��)�͐ݐ��J��	ݍ�`�;��w�L><2"��^��H�,�t�mE#g���8�2B�drz�|��R��-軏�` Qm0�)\v�}fFj��}9Bh:�2u���^���`���_�@��ݧ+����g����Se�-����b�����?u&tGJ���
Q��O�1���L���:wH����"p��c@Pv�4���h� ��R���0��J��f�8����d��y��l�(��t�f��@nܤ�V��R˕���6_t�4���eq��i�Y��1�����
����#��m�L����&�0�iI �2�
�d7��LW�i�;����\��g� (�e]���J.��Q��I�z$�Ae""�e�"y���@ �]H{���F7ӵ��X�k�-���c��v/g@��fw8F�Q����9��M���[�E�Zj0CSa� ��!}�9��;���J/�Zo�x剁.۲��T_ ��������#�ư�!�$�`<��_5�Ņ~�N�c���gU��Mހ�W��Rx�')ͬ6�!�-����SAjf���Pt4 ���UrNtOs��3f��-gNt
�����)�,�/+�`0��z@�Ow��m��@�-u�Q���Hو��uzۯ��:xc�^"�Ý�5�[ {sU��GKA�A��ܙ�(����8��M3�V�а��o�>aM�S�p��n(oˉ���ƚOR<-7�t����{)>|��9n�4�ZoR����tZ��g�z�g4\CS�&e�"���a�}{D��������%��A�)+� �p�V�8ǎ�{��7��P�0�<b��X�|܎� �uf�V&�4("��`��j|7���G�k�� P�nm�4��فc S��$�y��9�x�PW��lqc.2h6)3��D���@c��ҵ�K�{�A���EH�����?�)�U�G��5�N������b��z�2����ơ1X���2�?-+I'�}��d�S��m���/.Z$@Q<h�%�p7�޸b*Cl�5��a��i����n�Ė� 9͑�G0!�5��oĝ�A�<�U�Ѕׯ��u�80��V���%�����pĬ��Y�ç�����Q�o�	GC��5u���@v�G�Zab��'r��d��!��W1�����g"�#$�$��М63��� ��J�W'v'�D�xs�	a�G��(�u��Y���H���A�Zg?�K.QY�Q�C�R1��k�q�foa`��>�n������%lZ���o*X��n��FG��GVr�,~����L�vԛ�k�nט_�<��az#�7��N/�<��Grҷ��N_�q��*�ƿEO�k-����$# ����T�����C�.�.��@�k`f�w�!Vxv�zR���'����B��A|�<�98�wi�.6I@E������:�)�4*�2���M�8~���u�x�M#*�`5�A �5��o�ĘY�6���7ތ�+��+�>�t��$���a �{�Hؕηa�~�a$:~��^���4Hy�*"��s?�X�	���Hޔ��+"A\���`[���jO�:�*V�]�D_܏3����c���A�;��v�	 N^dP}#����R��v��=;��b�S��Ֆ�5_���eS��V&�����l��|�R�r�0�����i�/%�e	k>&_f�P�N�Q~��W�����B�F������A¹.LC�� X�6!�PT�ԥ���ϊ��8�����z�2�͆T�`���'�z^�"042�2��ܳq���y����;l�j�_��K(2�+!y#J�_���h��c��I� �r25vCV/�W��i���9~����ZA����� ]��n��ưU���hx�`̵@k-BSq����#}�f~_O3�����4XD%��Hʗ����cI�㦪���c����������/���k	��q�U�2M^�V.m��iLf�%�jA�>ߦ����uR%x�mQ�R��^p�(VI�Ia���Ưt ����]���Mg����aI��kQNE��,?"
|n�ċk�6��kם?���i��U;2n��Tհ���iE��:�'{�+4��N���P��"��<xxQ\by×7�h��CS9e��z�'/�M�lͰ��36ŀp�(�>C��<�mgw�Z�)ZF��4<��a)�UR��?!G�kj��`љ�f����O�2%�R@�HW�@Z�����b�_���:�-��o�Zq/�MSw?^2�Y�n�����P(Q! r7�2�z�f�`sS��sRU��&ĳ��� ��������Vl�n��yeg�J�ޘ�R|��X!Yʡ;g�
��r������.R��i�d$�L���%�d&��%tG�p����yo�*� �-	ǟ#��6o��s���2���!{ѕ�=���т���<oX+K�7��FW$��=v�\�92��^{�����̕��Sp�ѿ��-�J�2�k��Gb,{�@G�=Nܸ����#�����>X?
\q�z��O-��+m�H���b]zE����I��>@֦��S��f�K�#t��h�u?.Nݳڝ��ͣb����,�.t�5�3K�XuY�ɍ/�]�Y\�BTCN��QN��$F]ge�w3W�չчYf��1� �2!����i��s��� �{��9���.u~�yn�cwJ��,ӹ���i3~�:��K��j;��������Y0u����_�jB��}Y��<��&[P�^R<����[�+=*����Ы�W�/����T�2�6._�a�֪���6Ѳ�J���y*�O-����k�Q_�Ǧ�u'V���H��x
��1un�b��Q�����M%䖚5e�l~u��|$�Ha���N�n{�uz%��'�g��ź>#��|˫���C�����z%$��>�+��%GH0��Ц+i��·�UQ��_�|H� ���m��,�8ǥ�**�Y"��;�VA��ri��b �N���T
 S�wT��������vt�ݭ�NH5J^�P��P��0�m؍s���>���������59Q��ښv�R䞺g�kT���"�G��j�,9���-<s@�G\Z<�y��y�4��G[�5~�0U� �R�!�;^س���)(����i�HG~�cz�����"���1Jq�!Q6Зꄈ'X�A)�S�:�c�Z���2�����!ʪ�2�A�C����aS�zc:8��Z�b�Y���W2GBXY�h��Q�O��U&�j$�N�T[.K;��h4�Ѫ�T�*�Drseo����|������"N�:۾�%���]�LU��Q��e
ڐ�������w]�����d�0����K<���.��E��������]�\-_䊐D�_���Aog��3J���Aqh���!�Oc��S&��R�^pn?/l_8G�t�qG���h���M)5�5C=�>[!�������b���y��E�S!8�ː����}�(!	����p�����5��8'��iA��˳�)Tݶ�%�'�ҫB�����ao�1�؃l�	���9z-����F$���	y�-��^y�F����Id`�P>h���������&-CB ��G}�S�aѥUY֏�UCLUS��v h��bfݵ/{���1$��m�쿌]b�����N_&��I7�ESH�s���R��<8�#ώ��/��:}G���"����[0�i�e���U`dL�DR���p�r5{�B����H��ajV����\w�(
�{ҩ6���x�>7J	��.<o��~?r��l��~�B��YbO~I���1��jJwt͚�i��s��~&��!��J�� 7��Aɺ�l��<��F���{�2R��;5�*���|���!%ce��oeU���'�9yg)�`��J���CVߌJ+@!�X�/`�G8%
��f���ǌ{_h�+�Tsq=L�И~�*���NT��r���
:P��b���*c�?�}`���4���	J�7y`b5���v5r2@3�h:;Y��e �z�U�o}�����QmU��yz��/f�V�0Sf�m<~��W���������t\վ��#�Q��;��������`��CTE��/��\P���(�~?
�t8�l����硴�հ���U;3�]d.��L�z��,I��~�/�A�^D~���p�c���/��RQ���c]����ٵ�� ����+v���RIYe=L�I�ܽ'3���~�?
�rgR)q���lI
*q���(g5��6�m�/,�p�
q���0ifz$�I��S�cn�r�1(�\2s�Y���*/����z9��oMW�]�`O��rL�O�$��u���4�%h����U��O��ɵ�F@K��Lv�4
���8x���L��B"N��&��.�K��M��||���9��.Vp�a��[ofLG��Nh/l]�_nJ� �)ܠ<�i���#C-�Ӂ^ţg��a5��.�u��sTc��/D$9�i���o��L�BJ�-��Hy&���1��Lu+�,�ʟhg�U��0[���A��������w����@8uЄGay��H&>P�����l0����2�.�s�Ԣ�+ɕ���_��O���2Â��!F�x!��{A�I��e����N�cD\ 5��CF}@JLhr�D�����!U���륅*������{����y1�p@7��n�R|���:)n�%��}o�&v�D�� )���w{X��#�Y'C�<E�z�ɠ�:��Y�ҭ���P?�&�f�(��3û�Y����8^À��^um��g.~�9FW���}/h�MD�t��N����*�L��ӗ�P�
[<��c���\H[vW�/�/ 4���>�ɨ�u��}�gGk��߹k_��ҵ����!M����Ê����$*ZJ�f��/��^u��Y�\�ܓ����3xh�r"���r�+ɬM�}f�?�'��H��z��Q�,]�Nd�*?��v�&���o�_x/�Z�.u
��NTe9�2��Z3�w�3�aX�j���<��U��0��Ś�Y?p��<����\xR?D�g]܈��.I����g���K��,I>ۭ6뉔Tq��(�SL��$i��"@��J��ȸ��$�x`s�-}�&��Fiz٣������k�yT�٤��{a/V�V�ǆGU�qE8��q�Ζ�9c�pl<}g4���93^�9.ǩ� �D?^	���+��zh�#;�;_�ln7�h9&2��Y��?�ƱީTɻ�'%M��D�eKmxb�^B�r7ǆ5>���
��	o��Ԑ9�{�亩vT�@�S[��x|�z�<��#A�o���A��Us[�Hb~=�������,���&��&�K���4*�u�u	+�ntNc�Zu�wďUX]_b?8ُ$��N$�۠��M��쏧Po()�4�[��$Y�BT����Lհ�:CEhT��ꓲ	E[���1>����ޮ���W�y�by"F�O�A+8��bIΌ�;����u�,x0��ۗ���L��!��?[�E�a��XoA�Ӗ,�QaRZ�V@q��f�UWZ����%���v�����&��<2��M�I�T���	��H�`�o�x�1DhA�.�"�p�
i��TG]���ҡg��a��e��C�2Ks���p0�M���a�4h�����>6���BTv:���g�-mxj(j�9�BS��{�x�Ӓy"-���ײ9�#�9%����t�
�in���z����XE�"w׋�k,W�s)�`4�B�r���Ҵ$׆�y�|U�ʑ���S� ���[��3�ӻ��`�6;��\�CK��̹���oVu&�;�:3͸�6
d��X>��q\�qsl`�P{Qj���ŗ���dY���@'�c���A�gD�/�C�j�7U��!�_+k�Id6g�6բ��ܩ��y�@�M�mf�	���m�����^ɎI���Է�F�Ї�U��=18�Y��/���ϓ�S� ��uu��~�Ѹ�@��6���	���\��CoX�wI�xh����_�"�y�܌����[���ȨrB7�[齮�g]����N�N�:�Y��Svw�.b�3���E*vz���ov���?@��6��*bI&"7�,g՜֚t�]�)tc��?�T�Z�ĺD�$<�T�<�Z�h�����'?5�4�M(!�I�r���$�y�X�> &��sE� ��vP�[���G��α] �n9�tŬ���
�Rt���Ws��4����W���n���Ia�#}`/B�N���b�i��6���Z�,�xǾ*.��
��v�䗆_	�mb��Cy��>�b����︘�<�w�$�>3�i �'��Sx���~#5tp/�G(>{�zNWH؝[��r L>��=˄�aŦ�x&���-�ϣ�g��J;�m�|�=مGVvg�H/M�Z��n}mT�����Q�lj�&7�~�G��[D�P��Σ��$7+���8��/��"�u�bg$(��y�U��m�t���a��X_Lh��/�5����;i�7���ށsBd<��~���NWv� p���f��ō�:�_w[�B�	�Z���_�j�V7��Rܺ�9�(���ɭ��n15V+��L� ��+�Wv��>����n^�ɌU�SVУmF���'��Քԇ��f���~�RJ�S�x�{t��q��@����LE.��=��~.	�S��ؒ_�o{��;�=n��a��r!����է�Ǉ�^��C��{��1��	�BբB��΅��e�.����}J*qǫ ,������TF�b�����{"	��Hhe���6aD�ڢ����&����<�6�˱�ׅ�=�����R��z��� �Q�w��#�n������<c�`�R��4��:7_=�5 �<3�p�e�s�0�6�w$֐5 㨮7
_��*��W�e��앃�%�ڭ8oyb]��0�8�ըz�5�_.`V�R)2Ğ1�(�6���A^�s;�`�X�L�����}Q�<\�7I�Pξ�Q����*��D��Z���~�h�$v��{F����Yt�{��Z���6p��:��ڍ��	��g�ٌja�t����R���Ũ�2|���f��<��]f{v�Hq�♞\����N��ͅ�*c�O�����]�:���W���P	�et��d�a-�aΫ>�`y}۸"�!��j�<"��$�@��u*��3ĄO�	j�Xk�N�f���.�=b����7��P��0�R�F����~h���N��3HS$���vϠNF/T�y���o�Cx�땵0}q?Px[��T}`� �03<*{Ӳ�>慗]SxX�y��C�þ
!?��`��<��&j%�I�yT�3������Xל�V��ǲ��T4��}��gn�x�J ��Ɖ��s�r����Z��*=��w�Vv��`������0���-nMP�G�Eާc��f�F��멥%�*���2tJ�H+��beJ�1�'�������Rr���oz�Ew��(u;D�REh@+V#�At�A`�u�q�WF�}��l@rz��ӄ�{6d$Nn�}�_�_<SM������Dk��w��6$,J�{{zر��u1��(�6�jY�8ht�,�|�S�v+�f�)�8E�ErϧTa�.tp�[�E����;J�@��b@�pod`s�>���kӃK�$S�PC��a�q�O��	J�����nk�� �����/�?@G�?L�^��莿���|��Voa1��3'� �t�xS3�+�M-_�qO��}r�4*�<h��!Y� �.|�}��w�#��dG�ܽ�}0|�9cL9�aº �ךxڹ���:�i�F��b�W�;Pd	�P�A��O5���]~L���x2F������n]S>�|9FVV�A�|�NwSvn�`�t[����`��~ ��pj�U�����N���M�����<�#����OY��@�Ml��&����gpb��*�g�c�.h�N#����ǲ���j���!C=IiI�
���N��q{�O�w���=(�$qds;4nZFe4}t�'�N����K���3�9�5�*�=j��Y��R�W�s�����;(�����񡗫ot���4qn�^�号���e�W�"���T��zdM�,�a�
՞�Xl���Λ#��jI�(��K�g{��1]Ě�B�U�`ɀ�e|��`��9�l��>?��7�ꐰ�Y�e�M�u�{��D���s���u�G#F�C�����і�_�Z"A��~��Kݹc�T��l�8)0Zm����������ݳ+�y��@6~"c��Z�\���L��)�Ʀ��٣	/9�y��ݘ��bR�݉z�g�I3(L�&ϩ5vHM�}�w̴T����)E�fq���J���v9����Z�U
�͵魌����7�O�j���$�`�^�T�8-�D9�8��qN|�5�j�\���6=�1�#�0`2�N�|jo�ԧW�?r�C�ޕv曢�,��~�k�Wv��t3n��Xq�
�O���)y��IB����ѯ|Ds�d����G%�pOt���L��'� ��"�?<8��G��%�5�	�����9�Ys{�$kOɾ���kAT�,���uP����Hv A��v�[��#Qt" G�m���gh���JEa��-�H ����k��pyL��?����O
��>���x�R����!�Nq�b�sK��x�qǦʳf�����{GV�"����L��Cv�ӂg�?�Q�Eg��aG6K�P�Slֲ$�'�y ��=��j�pr�>^���� ��K�eMZ��(���=�H��;�n_�0��ul���L�ɿ���de�y�.!Ծ�l~��,ӭ��&�7�5���biR|�UF�D�x/d�Ek�"M��"�qv�e��+��73��m_
�������{�OT��~����5M�C�6�/E����А��-�9�IѾb�����
}�1��#i�����Ŷ����y���;k_a�$��)���AŅ��-���X�j"
���/�#�m�I�D�sK�E�E�X��ɷG(�S�]x�|~ٗհPY&�0������[����3�4���]�ŕ�Z���a������������x`b�Xf��KF��w�_�^�G���GU�_��?D`��ُ�F���M�y��i�B��m �uqa��x���L_�\\�c��IB����fo�\������NUHy�>�#yN��W���e�Ճ��pQ��.-����8�^3��X���7�pհ��i���G��]��l6�.�2L��z���BX��Ԥ��y����������-�B����H!�<�SN-��\�3��\��+$��f
p�He=�M	(:J�ϓ3��Cc5~�y>I}����G�3\������)*X�wS\���(��N���^x��~�K�ZUJ��X<�;!��|�C�9t�t8�7X�<��2���|���fo�Qo.��b�b�w�o���[��\Ҭ�?RU��%��}ׁ"�ҏ2j��FƲ��6a3���x�ݶ{I��R�s��_l7z�m(D�]G���4�4*�:�nP�
��|�dz�.Cq�����gn�m搪9eI�+��E�6b�y�{p�~~�A��so����V��$�hU�8�������L�e~,�ƸS�w��/[������E59���}�<�K�2*�(/�5�W��Z8�Rg��Te(�#I�o�s�������vw֖�m�|X�L.�_e����KLA�o��3_���6������[�K]3�D+���o[���Q�O��S�M(:�I-H�6�o�lY�տ\��'�:(����~����8$�6B��z�D��f=�.a;��3�b��!�ѫY�-n�H�����3�Mĉ�N�1]A��{d�u�� �����?2�C�n_Pr�R:Us�7���M$r{O �P�u0*��4�ʈ�n�2d��-���tgl#�uڞ~���Z�v2�6����G|�G�Iv'O~b�ha %�*I�iS�d� �7�7^�إ�D�?����L�ɼ~�b�>[{p(�0@j1�2Z�m���l�Ѓ�IU^��[o�ߐ! W9���J$B��K9QR>��ұ'�uR�AJGb濋�I��ϧ`��Y��n��kBЙ?�WH����0懄�4O�!��3�OT���'�}( ��+��=?��8�"�,��Y&��Ƴ!\;�]�>S/x[��R��k	���ESY��wi]���j婖#{?r|N���*�\J����|�?'�ߔ���y��v��J�@�u�R�8��Q�u���cy���rknc�h8�f]$��c� ��9��C����;��K�>����2Vڶ_I�dd�mm�0bfA-pgڧ�W["5�G�tE�\QYM�,�_��4���x~����2v�C�G��,����ڂ'���G��#�m@8�r�L$o㗌?b	�11+�_Y�(J1�i{)�6'��k��J�,��#�Q�����Alj�2�e�����)�8G_-�ߢn�ȋ| ��s�<��c5� �{E���VH��Ȝ@5� cU��A�<k/ߏ���U���/���,%v����HXK���ku+�:�&BJ9"��8���5��?��l���V�4�hшAGn7�|�P��c��\^W���UWMb1 �)H��C��w�O���̃�T2�r�.�rCi7���x�L,��_5gF4�aԳ��S�0V����B�5�i���w�ה�<���M
3�������C� ����a�q8��<#�i�L�H����qQ y�x���t7���f�R~HUЃ��}�o"�6�~�b��m"1wm �q��o�������:��JZ�BU��;b�P��li�(�W)�\����+�ǰg�������
 ШgH4��� [�A��8tl��p+������e��8
P�c�YE��(�Pl�uH�TTW[�]��1�骭��d��fa��R���͞1a�@�!ʸ�����Q lν��6*�l��c�0�L!,T�"�|W�_^�C�(�9AĘ��$x�\�2{LWӅm�Q[��{>���.r��IS�{['����h�kF݂8*�?W-���⡆9���g�	*wq8�}�t��پ��Z�˗�P�A
VD��+e�^V��O7�L��.l�̉<U��G��V)��N���f_��j���Y�a�Í��|�&q��2<J�$VQ�o�5��(/�l�&Mo���C���o.��Ct��g7����F$xXb�����׼�܍�	7��Ye�'��G�IQֹ��Y˯P���F�A,Tр�R�n�an�$hrʇ���+BBg��; ��K��;b-4#W�Po<�e���'JcZ��Z�Y)�L�/f�����b��G?~3��W����՝�L�w�<y�"�Ǭg�����<��İ�2�on�!�-|�K*�������d��A��s�b���%�{Z~���Cv��O\����Qb��t���pS�4�y
�z]2��|6u�%���<\|�I�67d�^lo=Q��w�o�R�S~@f4׍��$r�㼔T�o{Ю^��
V\T��� �CԤ|,-`�!����~�|l% z�C3�ɋ� ��4�K:�5{���Mk�k���d���~���'z��w;j��&&����	4<>��
��~Y^�wi7I��'9��.��O}�����AMZd~O"����}@H��B3�R? �W�?��R�����;���H���w0�Wz�T�z�#���� �Qm��x�4�B|m!�rK���BŽ�3H3�Ի��R	_�2^	�O_5O���m�R1@� ����ǊV��g5r�Դ�0�n:cL~��n��?�<D*��Я�Ki�*4{x�v:z[{�Q����IV���:R��A6`�S�0"M����Jq& �N)u;�_��|���Bh���6�O:`����iLIψ����y7c�\�}�����j� ���xy��lH׎��;U:��O��D��)u�2�a}m�녱�0���)n��9�4:q߆�>�p���ŝ��ߠ����/d�b��Z���d� �g%;�f��n�:\��n�Z��5�V��I9 �X�\ʘ�k�����Oc5������{���m���A�^�%��=������uP�'ȹ
q>�����}�M>Ol�|Pj9�!����r _�T�w��Aګ�#�yb6�5�J��c$��U�R.��[��~����Ŷa��i�W+Ѝ�-6���,�74�����Z|4��ʙ:�/؂~����(�7Y��Zs���σw$M�"�:	I��Ԋ�P.͹�Jz��M��w��ĆN %����#�,L��7\�0o�`t�-f��V�+h"B�9ԙ��wS����pJ��c
`}�wO
�?|2�a��Dg}������ڝ�䪦,�W����ȧ�;�#!�A�L=��c�=�nx ���4�P�<-�݂y�Օ��t�)����M�m:��J��Ve�i3U��Ew�Y��wBc����|I��٤��(DMy<���6A�\��hJ�����yu���aT� ��n=�B����O6�N����do�,����u}n�Qy.I��feFm͔�Ӱx�����T�_2�Z[R(�Il	r��*�D��=�Q�q:��1=�<k��!�%ݚ�(�H��m���<0��ș�cӗ2c��'�pv�A��X��˾�f�n4�O�����)4
o��!�J��~PE/Y]���Լv�[>�x2W*�<U\? Q�������6i� ���)|PqnP�r\gK��F�C�r�c�	�4x�R'-�� �>dE�x\�U���qo����]�[������}i�V8YW6�a�^������C���|Y^������U"��scƛ�1�D��/z�
�iwM���-�QS��g	�샌�*�{zr'���ܓ-��ktxW��Y�5�&�j;5a�fn6�%)��	Uew�7���Ǒ!�0��y�N�|��'?jr��g����*3��
'@����h���+R������mD�񅔙lsRP�{A48�����N����ٙ*o��6�v3�1�$O�4��,�f�G2-Q�K�Ӌ�[4Ka�ay�FfYP}= [����n�K��_ >��z���΁�N�)#[� ,ݏ�@$?�y�V����^ֆ퀠+1<�H��&�l�]jԮ�B6TY����$�4yPȣ��	��$�&w�iѝ�y���s��zznSX�E�y����#,�KPI�}���c����b�6��0����J���K�vmL�݇���1n��tO����63���v73Kl� '��n���rg�'�Jl���t����%_v�HR`��L��A�3�c$�ItN:���&���<��>/HY,�淹n���np�h��W���kK�B鿪M�5S��{B���ȑU̓�������g���[�	K�h�`k��t�f�J�FTg��No����)V���g9��=�����U����q����~�8Ou�t`��'|���������]Q��T�^H�����3��,�9kм��E{��h�����=�AmrqF6&�TX�Aw"N/a���<���!�� ح� ����hVg}���^8��Ree��� �P��
r/N]�M�n�^�\]�l?�`���)���i���9�3x	�<�;�Ɛ�B��&Y�P* ���_j�&VՇ��D����R��dW%�
?���ʲ�>,��d:�ò�	To0��N�^8%�h�xF���_W9�=Zo	;I[��6��m*��v���}�����c(��;[���Y9܁�d.�Y~�=�t[��O�b��7�>�k�k�o�l!�8�P�練�k_����媸1,��k$�6~w]����Y��7H��������S�����o�0U�ƆG ��OCu��I���O`	�ʙnǾE�I;p~D��h�|0)��`�p ����r#1жt�N ���<L	̯���ݺyw�徧���G�lT����}�u�Iy�<S~g ��g�1i)O'��9�������]Or�B�S1�5��PE�f�|#M���)��gqO!�q|���03U��f/B����U��&��?`#�������>�5��$t74����0ڴOY�7]�T�8 �g�v��;�Cg���B�풠9f�#�7�mSHȂd�je ����Ζ�O�E�j�S����������^�h�E{�����l^�tu�ڡ�q �{\�1FP�Rzk���"�?��|Z�T[�'ے]l8I��eSLm<�a����̹k�*j�q� 7�Tߋ?��&�aʆ 7��fէJ�D5��������s n�W*�S��@'������S�J����� -���M�qɚ-��-��b��x۲7�$�UC��Q��LüY�Ù�:�x�Ϭ�{�	m�����GL^�����őS���2|� ��W6���^���v�O��J���	��{x-=������9̊0�|o�ېR��$UU�y�8Z��yK�*˂W��3׳}fN��VKr�m�_��l�DyjtNc�"݋x���5�(#L�	~	D�k:2Jz~������O�8��EA�/2/ |)8|_�)��'�(�.F����l� u�#���EP�Qɯ�ۙ%���W�M��k _+�de�Fl���;a��v".��mRl3`Z,�t���:���>W��s*D��>eqm�*u��pO���csF�|�[���/~��O�k��S���	.lB^�$�5�6" �sAƗ{M����������N�9�5�q�k�|2����^�|�%c��*y����fL��Ȗ�%��`��B~ (�z%
� ��/��������&����IÿlS����"x�,rDq8V
��`!�	����2����`ĝ|�\�͂ނ��6������zp��{��UY��k�zJ+�Z"N�����ĻR����s@�?o� ��=�ֻt�J�H�z���u|Qb��fX�Q�*�#a�*�	{���Ϥ҃`0� �h9C0����aY��� ��r��f�Ѧ���T�����%B�\h|����2���6�+�<��r�sremI�^�W�{��UV��d&�M�5�0N�ݛȭ1;٩��1���P6��n`\�rt���Y���j>+�Wfu���CZ1������B�+��+dxr������o��k1�B;�(������8g{P�[ü�Z�/���ʫ�+����+	��W����� Hb��P���2�����=���?Z���w�_�Dz�$ģ~λGp�̖f��e8�`W�y�e�V�kJg�����21 �@H]�n_0`��Mɀ��Tr5Vdm�1�F�[��-��7�?�����o�M"&���S`��I���V;�Ö�rEi�',vXt0�������4P<���n4,���ӷ-�	SE�1Y 5]���O[P�E�IH�̝�.���oaB����X�	�Rh�S�����c�p�3jz��6���)SZ�"�'��NuƴꊟH��Uæ��A�F�P)�\u�_�Rn^��4���%�ݧfq���f31'��2��e�xr+.n���8��Z=�x�/�W��ކ���E�NJ�x�����C�<%�nb�ԏ�w�D�ȉ�B�ۛU�����w}*��m��Z���蔶�w����L���.�W������oL�&�(7-��Z?ɫ	]ke�1[m-c�	�=�0�(L��R�G���
A��Y�C��Fp7���c�x���Lkv��X�,{���@�Z80w:\��9��6���z_7�����*q ���Jj[`�^L�U�]��|.X�7gj~�Z����"��%�:	G�����.3����Ӷ��7674V�K]�Vt��w���X���b0ûV��� Ǿ�]���b��ߨE���֑�U�sc�'P�PR�.�/)���>j&�����9�)u��V��v�5ra�� ��Z���F���cH�[�~�G�ueԁ�A
������#�"
���	�ǁ{+M(�����O��N/��+1^�pz�h�?9Jˍ�?�dlk�;H�i��-|�(*�`1����F;��Ff&�b3���z�v����<�=u0 �R���o_�t���uE��؅�&� k�W�j�F�,B����}:V�.��[:v����Pxz��iI7�
X��N7G�c�?r����J
��*gXMMǿMT��o��n����b��r��BA���W���7��\�J.&����~K�A���̢�+�y
��dj6��.ӧ� �����N������h�#��{K�ѭ-ѩ$�7�'�ɒd�.z��j��)a��1��b�kW�-�������p����y·\�7EXП��6H��>�w��˾��6������p7��Vۘ�tu�4ۗ�<�6B[@I�XR�'�T��H�[~� ���~��ªn�	��]�OZ�J���3����P7�v�Bq ���Т��O�d������2,ݠ��M�D4���3 Ѻ�w�#$���u�{"{�Q���n!�Q6�>��㗇/K����C�W\CM9�|��/����ōF{�v�o�әяY7��\)���m������U��:��m�y�����VOW��2u���kl2AmTRG��dˈ=圼�/�D4y���s���)�G��gO9Rj�q���0c}�H����|�-�@�=Ǿ��^G��p
k��^
��-�\CQ*�qŌ��ŊbGk�휏4�M�(/DL�w��?Ęs.�N�PL��ݯN���DyiJ�{�B�e#$*_�fCs`��[嬅���k�$�p(�!��a�..�?K��4湑'�������������3"_p6U����i��=P2I�)��5Y;aX��e���0Igq��p�uW�182�T-�J�kpc�X��uK��;�P+=Wİ�?���'�f�>�`=�>� O�/6�n���]�|��;��ʁ6������j������ b��0j�Ҟ��ڟG���fS8љ��ȝnc���H)�ҽ�r���_u1<���co����=��@R������c�7<�9Y��k��rV-����T��($�ǒ���&�l�L"�M<��\�'"��'ʘ�=����3"��ĄM�7�;��?%��|E�bH�t%5�í�fF��8L=V�B�Ǐ_^L�1n�]�*�x�&b����U쏖l��j�\�j�E�O��I�d�戺f�,;̅��81�l�'���C�9�?��Q�0a'��0o�������Ͼ��9SD�g�:������R��`��d���9#{O�����y"��޻�M���s�J�hl������[�c���bO=o��;�#o��g�!x$}���;z�w�ɂ��:��_m���o�#��z�\$WA�8&���E&��`	��pD���شi%mۖv��:+K�.�R3�/���Jc7}�;8H�o�w^�5&?x�.Πvl;5f��P�y�>���t�Ӣe�A8TLHP������w��p#�DS���<����_��ű�~�L�BZ��W�C�f�����?�h
�k ̐E���u���//a:6�Zٙ�-��R�f_m�[bu/��e�1���i]�fA��� ����^�@Q�>�,�JV��i>}�.)$�O�Q�ϸ��ĞK	il���kl�m�H�������
 �!q5�j��H�qZ�J������y�уJ��Far���>�r�����h�*�RS�U���D,K;��Ϳ�:H��}⧏�+�^\`�>�-��@F�,�����$�Q��zK\L����U\��y`D�{��)�@��c8M���!A�Pa�3b�u'-n����H=�N�ƚl�{��=�kb,Ug���u�2_�4�o�zie�"��>:8�»�^p�GƷ�ġ�����*S���Ik܄�b����y���|$��Q�l���!4��Ma�7$:�!ԓ�7pg��O"�cY+Uz�\e��5*��vh8����ꩦ�c$�ڢ��Otyo�j;U����'4R� p��Q��Dקиy'C�1Z�h-�f�A��x����?�@�0ߜ�V	�|$G"��`{�'B&��C�������e�U������S(�)�� Oη��$�l���BXEv�3i��b�o`5Kv��Y|�\_��K��nJ�ے��r}<͗��?�L7� �i;�F�?a�$�V��ӥ3C���7:�-��S�NT�f�@I��v;#�i����L�|�����H�W��0���6�H� nMP^'2�A�"{�څX�߉1$�0jak	T�?9�?�#;(4���������krT�_z���z"��])��D1-�UMvR�]����� �¶Vl^z�a��T�������E�bSX)�[�4�OJg��ɒ���(0O�����w�V�<pz��fZ&3$����� ��޹��7�d5�1
_m�����'���������/nƴ�N|��ԯ����q��ηck��Vg|���}�!볔��3���Z�>�q�n������-�A�8��@<��0j�7n7�������&p_�Ѵ�є�	��"����mS
�s@7�o�ֵDu+��I��"�eN.=�6�OU�1� �˔�j��Jt�33^+�%�+^��|�
��G�+��B����p;4�G�]��}��/�KR̢#��g}f}��Eώ�w3N��[�n���W^wv��j������P�d�B�y��d��uԍ�ͺ��Z���k��z��EMm�k���3��U�>��8෧-I��M�r��(�2ދ��|wr�GXa��f���I�^����ן�2B<�hG�������F��Ӥ�/��!C��t1�o����@ꯂ�n)��,61gB�"_�:�pժ'��G,E��)�?�'߆e�0Z7��un�G�Tch�����ϐz$'���J��|R�Y��q�����O�K0Z�qG�!���l�����e�����swf V@�Ǧ�͘Kw�p���%�σ�&��ؓ�7Zj�:��jQIz���5�����syAc�
ts�����l(�V��"G�1ƌ;5�Z����J��PU嵄�y�y?����I�Yꇜ:Ռǥ��|���1��[�<+v�����z��6��wB����[�KA٨��Ie��~�U9k4��jk�G�^��rpL����F{�ʘ�7ͪ����cm0caC0����p����F�v-4��U��;���v�����	M`�4ǥ�W���>�W2t/���%Uwc��n��R�J7p
T����hBg���vz9m�r�r���o�eC;����lz �f��X���yƁ}����=�>ֱ�b�	\I>����.W3�=I�
�-bY��;�>�J	b	����<.�����	��gs�]�XC>ַ��%C�qR;߅%ڇ��D*�(��Z)�M㥱��]��_cntT��/h��J]�#�JA�LRiϢ���jgYQB�#�,�#� �TƱY8^T&�G��6��}��cߡ(�o�W������>+�  k��X�c��� ~vdV����_�sؒ�Ldd�	C�����.x�b�_B��pzk.�;x�����j���D.�!�g׻�i�ި>��Hޖ�N��R��!o s���Fx1���y�+B`� 'A>�Q��\�(�v�?�I��?w�t���)%UApd� >��o���r=��i�� M�kG�'�י�Iܗ�z��mi�%�:�6���(��H�xE#���S���x�t���cv��m�����lN*I����T��p�g��Ջ�앙^
^�k9Mk.�T�y���X1p�#l.�#�� ����@>�#���slHJj���%ho�ZV���� ��a�aju�I�An1g��F� �֒qw-���$��`�V�S��U�ݒ�J�ɽ#�r�=;��i!E��^�x���4ZDP�2(�x��݌s�~Y�)��[<�f���g6^�)�q+[g[�z����n���c�h/������Nb���V�b �r:��
Vw���:�p���o�ǐ`�sg�W#\{F'��,i��m5*H� �,�O��]u�i�~� �nTH�T���(��	q��fh��1
%#ܱ>>I��hRvNuTq}�`Vi�Lp��nzVK��p��dʖ�:�PI�ŧq	2�Xx�;���=�cnE����/�q�"'��M ;��e�S�5e0f�dCy��z��L?�K���QK/�h�h���;�?,�bHJ�����^$�^�_T1���2:sg�S�)��C����^96n<�:���L��*q��礗�^I�Q��|��NR}�on��H�Q�4c�Gl��g� k���K����[��AT3�/�A8F�4Џ���z6 ��}�N�X�+��a�D������֟�>���cp���E�-7��hs���g���}�8�5��%�{�͖���qV�0���r�ITI�!��m�Q��^ U�B_��K�8]��E�K7:�f�����W�19p�н���}w�X�E���W���?8v���qK蕙�IQ5�����@�(C$W��8�Ȼ@��m�χ�$��o�1���1��/c�K�b���ߪU�'纺�ٻ����pJ'cb�L�u
I�:CD5�1�sN,�ŧ{�h�ꧨ[���+�,���Q@c�;�����m ������[c���؛[��# !ir����T�"B���n]$�2�P�6
�Z[jH�{9j�"�yEwN�}�gɔ�P(��n�b�s��i��c�D���6V�(G(,[�?f�p�a����	=�@����\���rL`�#z�)/�{5P����;�Ң���R� ��{�(.�F��q��IFrc6�;!�63SB��ȿuCsB"��@@6�e�T����	e&�ǯ5y͏Q��#���E{�@��/���wsYY�#��L�x9�F����G� ī��	���w�;@4ݍ��N	$U��Z�.���tM���Ы=����ֽs�c0n���q�I�_Q��y��+���RXTԖ:{��4�H�Y�\?٥�Y)����r���r*�=�֘�&��� ّU�$0z�TD��k�4��4%�)�%�Pc%,���9JAMS�Ө����u<[��\�p)ϱRn�Gx�C2���|e��3��r9�s�b1j
R0����U* [����Xtc�<R+L����4��Mw��6����xr�|�˾�0��iѽ�8[���4����>A5�ܰ�6�G��g�o����"�A���T
H�)e������lm�7���籂q�.<�	e��_�'�r�` �������*���O0#���RmɄ^�-��nN^�73�.z��H��ޕ;��	�ȯ f]~��Q'��[��zҳ�{�Q�X�eA��[T�E�n	Fp��[�`�F-��Ry�)�vmٓ�EM��K|f��a��O��@��L!���P�pJ=���E.ֲ1 Xx���ɕ�9x�q���X�Go��8�R��O�>��Y�U�-ⵓwþN��l�9����7Z�����$3&E��PS�ٓ���s��d�:/��{(4O��G�JB=6S�)�{�?K�A�˰^
v�[ٛǿ-M=�%cV�ÚR�� ���U�bU'O+-c^Eo�k���w{�L�Vy�TZa9��)<g�����Ļ(/E����զ��7������?���F��@=���#��qM\\�c~vM�o�;[�N)�y�k�2�ǀ%���ਯ��9:�Ι�}R�>Z[�?|�sf��\.��l�Rۏ��D�x13dx��� #�����l�;9_"d�P� |`��|��[�c5Y��	�xc%䐽��5AS�D�]'n��T�g��0����Tͱ땡Q�B ��N��@�?-�S�ٽey�x�Y}$ Ǚ7j�3|_�ao"Z־H
Q���S�RRZ.�I�L�ߦ|"bʢ�H�7u�L����z�)x��a]�ڔ2��6�}D�`�i5ʽ{Ưq�_����e��&k:������(���>���t�����E�ƌ��qJb���]q�˓�Q*�W�>c������=�oEKɳ�))<d�� Bd�ca�p�-ե�M���g!��K��=�'5/N����.�e�ȍ�k��1�o��l�$Tia���#:�((_n��c틼�`���_P>5uӉ�Z�d�s|�&�ԛ��Nh�S��jӽA�HQ.�:]�ɜ�ͺ���&���]���!6�[�u|�1l�~�� ���< `��Ao/1ކt�)r�G!!�''Co����ҚdK���=y
[f�����g���x�u��ES ��q���2���.z�p*4��WN1r���M�y(�E��g�;��vp�T���>�P����4A��q�E��na��|��ED�L���!_�C�3���,r4S�����	:���������n%��n3�}����kTϢu��Z�ڥ��6��-���r5P����^�Z����a|��f~�����'���)^D�a�p�I1���p��{%�z�RＪu�x9ĊM�4��%诠�a��+h�ڤ�@��;�}�#a��%<?�e�x��\�g�������MCՕ����Ԟ�ʸ]g��R2�l�Y�pl�]vȊ�-���Q>cW�dN���3�|H����	l"#4��Z�C���{������[�+�[�7B��>�7�[�!��;���Τ&�b$;�!2�[�m��B�u������������#�],�0\��]�wp�U�g�3�=��f�D�;jlŢ��Q0hf<���'��Y�
���[�|@v	�2��/"ߛo:i����^P��dĔ ��m����c�����()�v�e��]��'������^�ǵ!����+oz(ȓ�	R�j�^�ғFu�/@$�.�W��B1��&����N5�!K��W�����r-�2m��_�7�ûI�����o�D�~��������t��l�%�$�x���[�RV����z[߹
&x�wwy�)�uqO`���>���pdԷמ`N���Ԣg��>��m���DH�ɵ��D
!��-=eۜK<��fс����I��T����,���J� � ����X��4�$��`w�z�ّ��*�",�b�U��r�ӄ��a,ս�f��u��Yk`�T��̵=�y�x\.����$��d�T�!��I�H��~�V ���>gDTM*�>����A�P�OHK �B�v}g!��������+�
�I,��HEŨ��U[a{�[��5��6�>���b�<� ����� ��Y��hu�Bg=������[��M(`�"�%��O ,=���L�G%�e�����ʂ;�]\��Q��X@3���E�t�f��2��ch2��{��-A�O��х#tm��-3 J�o4 ny���uoGU���r��eS���Gf*�&_�>��,�\�ld�E�G�'��3h˂�ˀ��4��,Q�|�F��9��;�i��y��\ �c��'-ܥ��7��������s������~�_:a.n4�>��6�Y��s�X^"�����,�<'KF�a[��7W8�]G�WF+��=��ʕp���l�]��8�9�Q���@J�4���e"���I��8��Z>��UF@�.YF��B/�4+>q�A�����,ո֮�\��&2��+��?�%u|�����#�0�h箲�ƣ(ax~���F7�AP��fY@t�r��g��Dր�����`���C�U9�e�0I�%��x�a����,n�<�V �
��M_b�R��s��W�����v�5�'Gt0��0���n����x�dɗ� \�0zt�_6�%f�:ͪ����9��]SFJ�v�u�ٿC�C�������g,m�y���8L����moT$$�I	�'�ݰm����t+a��+����Ѣ)��z��Di�ST_	�9���l�ѝ_4�9F���8�ⱬ���K��<�|]�vCn'��c��&	��fH���KBec��O���m�r��H��������*`@#h��r�Kly��Z^Mt>E�^���;-��|G�C�1����c�V����)��@ÌjT'A�H��e���:J��$Cwa ⾘1#���Ej��k� �r	"�j�' ߲��R�Ἦ��$�4_��.P=$���������!X4���7���H��o_t��o&�`�ꗊZ�sCJY�4�
��nJ�b��+�xD��A���

�d���_��!lUAdS�ϰQ�ktS61� �����rɃI�����AhF��"���9���Y��m�\ۯ@��Pf(S�~����FA�� ���5YGz�#�&H���E��P����uM��8]�Leq å�SP���W!Ұhy�Z�K�Mc̶T�I��
�F�9��U��	�������ڴ��e��)N����~�Vx�\]�Ҵ�p署_���'e+��[�s��#��.�c�.�_����vZu�3/���{�z[�E�48����5�]P=����P"�������&�CN:�q��r؄&��8��b�Y����WK�g�<<�~����m[fST��jN�U�� S%~���p�@� 9h�o�^��Wɜ����6���?ʎ�8����!	(��HJ��~5">���4�Y��!@x{K	[�] ��^ BzU*�|`�wSU۔hIp^��b�E�����u޹ϴ�A�rJ�3*-r�F�>8�G��`��c������iD}�ve�=��E������Z�?kt7��(ϩ�c�A��ɞݠIr�V%u����*��� yi ��:����HyBS�{�O�T_06R	�`��~���Ǐ'�U;;�5ft�2υ�Yx�ylW�
������ �O����jcz�D]I65����"c�t@c`L�6l�IU�0M�|?KR���ų���Wk�*K.�QE|*f,RVsy)`(Dr�ȩm�p.������������GN!��&-�'�`��6;&,~|��0;��)oq���a`��/����r�ʝ*"������6�u޼����8��HQ���%�H	%���i�:{b���)&�"�9:ݏ���B���t��e
� ,�"�F ��w�c�C�m�.n��_�OɈ��b��������P����@�5cz
�0׸3�b�>7�}�4y#���l���D]fC��O�k_\a��:�1�x����M���"+����5U�P����d�-��d��ӕZ�(Xى�U��ƩӢ�O{{��Q����>{+ғLg>�^���ș��?y����U��%�|�%Ѐg?B~���UVD<�����oT�g����������E���#_������O���R��Ve��kPO�*�Ȟ늏-���"��@xo��&��c��Xxx�Ԭ�O�QzC�nc��Gf�S��F��s������a w� ���jd�FS��)����X(��T���j�=ې��:��7f����-U#��W�AS����f����ݤ�*i�.DL���4m8�>�YS֋��W��%���=a�[�U-( ��k��/��J{�BG��ɩ��r�+hU�}���z�O������)��G����	(l҉�_��l�5˩��Ǣj�n���2[#�BP��xL#b�ȸ�ļ*�n3���|���(�Ed9�ꠃ�ưs"���6���CU���A�@�0
�%5��K��۬i��S�mUƵ�#���7!Iz�re�[����W������yly��Q7���GE2&��3��v6@��aR��>_��e8㝋�c��Z�Q<k���������v- ���k2q�¸3���{�+1�z���y��]�2�h��t�I�����ݸ�̶�	�[�j$���`���"�B6q�������H��4��&�+�[�)�2W��I�A��X�Bꂫ+!`e:H��\T�Q����S�:v�9���"������	�k��+.�~T����C�y!������~	^6[�׺���z�h�Tkb`�Ӝ��-�N��Ɲ�8��-���N��/&3�g�اΣ�A���,��F���
G�<f�7l��/`��k������O�Q�6�$]^���}�=��eBI���ۈI	s:p�֭�ԡ�t���~y�� ̕�1F"b��@��:у�=� ֈ���3��[�Ѭ�k5��g�Dy��ڏ|�m�Y�c����7�+SU-Lq��@"�{˩���9�m����YY�����V	J(��mR����<n�o1mGe}�R���4�A_��2ծ��f���p��
G��6p����i�% �++˿��S�*����/��jb��H��E۪ou�R��^�_p$�܈��B���!W_�ֆq�q�0B�"n=���㨺1;Jd�-U�������_VPq�70�p���=��.�������\��R�-\�y'}�v���7�-�7�x��iO: e���\xi��5�c|cG=k2��B��C�8�z��H���E�:[����\5��eY�L���3t��d�Φ+��sOm�E�8��!r#�Cx"�q@������`ȹ���|<�t[]u��"�^���jW�@�\��mJ��Wi���fb˽y��޺*��!x4����|��\M��������ߵ��kSrYgW{I�D<'@��{6)��F��3i)5���l\K��9�1@��wT���RO4܃��Y�5Wp�T��|%��e���1�y�2B��o���V��H/�&�8@�"�̇����*���>wp����p9�]��	�^{u{'�Z��N̠Z\L���A1M�Kw��x$�X<ҲR�\�*���P�c#��2}Ɔa>�E,�������L.|B�Z��j+To���O�m�#�!�?МQ���'���O�!!I
���/��,������?rh��5� �?�����.d����
���wIqa�Jq�ӮF�E���S���$�#��W�`m�h�)E��īu� PKuT�O�rخ�����!&����9t\�?�S}���D.��h^�l�4s�*��� �i'�����fp�e�b�Ek�蠊���j��<cH;�|���@�һ5q0�M�I<%蓊5އ3 1oŠ�=�3H�yj&g��@ͰU�<���K����M�Z�^���{k���۞���&�X�~��J��_��-�.<H{ϧF�_���~���>(b�?0��¿΁�>�U������i�x���neX���$3Rl��x]c��ϢDʅ��J��|*}�ƨO=!C΀�1j�\��8��s�p�o[w��V�����r�j����>����u�Y�A�L'ڊ�|@�Q㒱4��� ���ի�j�\~ ^�lE������ɑ�%��C	,!ʈ�'�<�G`$iRo�.������&*=��g.�M��m�^�Q�w�:��O�{T��B֭=����1i����[�8}��P��͊^&prJʇ3š*�h҅e�CR�^����Uy�{GG���ʅq�c�.澆5$��\�@��T%�ͧú3�Y~/w}���1Φu��u� U�G��W�bטA�.�Z��R�`߁�T�j	��p�Y���4�,�}�Z8	��Ϡ�N���g�ʘ[r�R���'�Y�_&��#7�x���F���F��"��a�bk]��'���嬾�2�.Z��O�Sh��U�C7o���^Ek`�AxF�nO�4{*��VSR2R4��T��j7��o�N�9����^�CVP�ԯ���VO͖Z����I������-�I�5�7��)*0��_��U}��9P���Sʓ�aD/���B��^Ј�xT��	����WCU[-i��Pa�P�×MQb����T��gܮ�K�g熱�^�͟E��t'm#�.u����wZު��q>��f�h��q���<mۡ�(�GI��=�ӑs��릯�NۀٲOJv�2�'.�ky&� ��5������Gæ�t%߿uX�>J���> vo��Q�2���Q��[���>�i��$�`�W�֌��P!��-�V��L�]%��E���^��Ћ/ N��:�˕�Ƃ�)W��?y)��/����������ʋ��$��j���/X������Z�l.[Iɍ��}�}�ɶ�O�1�S<Ξ;:���&1�a�ɮ!E�}���3��)�*��l�Jd�L��U��>��6�?<G��Rɔ�8w{��1R��3���*|�� �E�g�7���M�����Q䮍B�������͑����+��C����K�}΃���>��1][����NO�֋0d&�����yip,k�Q�;�,�uOG?1!z����> �q���n�FK�2�����%���!�b��.��<�����{@/X�X�JfaR�7�y��{k�ۣ���ϛ�{�"���e|c�.�����Л�Y��1�BD��9|֊=�<{�M�!cğ�΍��HHn�.��a�N�J֘��I0�+�ɴ��f�������f�_%����{KdKP-`#��N�䥱�v�U'��#\����}k�1q ������?q�YCEvK΢���
��-�G��bgn3�9�G脕��=���z'��!Y�P\���z`���w� �� v�.p�p\�ύ�4�oɊ�������cx�)��j�����gy�j��r�W:�U�K�c\�%��<��_߾Wu����5�s���ݸ?x��g��)b��yH��9b�!S(�Y}���@�nJ3vޢGly`uS S�$0��[}.J��{�U#޹��=��?ɪ�Ec�D�2�v���f6c-�yl6J��;��t
��I��Wn[��A�U�_i�<�Dn�W.o:��gO�f��3�y��-!�{([��::z���U��w�~j/Ģ����0���Hi)�����Uz}!/q�B�i�b�-�Tڪ�9�~x�1)J �,)�o��I�E2����/wa��l_���D��0xb`�g6�򨙈��G =�/sGTf$��ʧ��Ɛ���~px-}� �no���T���E��MX��cKv��0��d�7�q,��X�bc��R�S�S���L ���(���b~| �jZ/D�{�q��5̶1sMb2��dy���&�]oE��)y�7���"5��+�G_J(XS:�/-r滎g�(�v/���?�<K�}yג�)��4>��R���)#�v���Wq�� �t�!�Q4����G����yO]����
ɾL���r����R����h���1Oe@i)�5�UK�{���s美�D��\��5VȺ�{�7b�O�8{��������e�1W� �6�,K��$��"��#>=^v��0�����G��+׽��	��ŒӄL���	VY<����JCy��H_����[��V�4���ؓ��4P#��i�Fg*l��l4�0>�_�]��uc�Ā�Np����Zk��z�ͬ��<D��reJ�r z��0<��A�Bpe瓏��,b7�}��v����j�Ax ]�����j����(�O�:��=E+�q#z1�o=�l՗>A��a���*�LMI�Gmv<�݇�.�����)�yћ�jl9���7�N8T�uu7)q�b/ED����~ g0��5�
�y��($����'�ZSIf	�	�5�T"���Ϣ���XnH�΄@B�mt�"�k���M�E#n��;��-X���483��I�%�m��,IJF�E�y@�N&y�E���&�.�(�U`¦''Űl鵂B����]�aee�T�.���F D,A���	>�ʑ@�U�)u]��쓥�mSoߢe���_��ײַ��[��[W �N������U�PR�!�?ALW���W�q˿Cm����th=�$�O�y�p��3�Ԗ^�CRɴ7X���R{8B���D�n�����.�0�LV7�(�/?��IX��{�����be4Ɖ{K���n8{a��-Wۨ>nO�ʦ�[�-��j:Jl�`��*��k��`ݷ�@Xܖ�,���?Ht���i��B�+�5���u�c�d��-6>&�!<���<��N  	~�s۠!�U��j}�3���%�-~��)³��/'ϥON�FM�(N��K9���v���ʥU��[���F�����uRUiI�f3�F���HLŊ:<��[6UOl�9�oi+H",���+�X��l�m�A�}ύ��7�.mދ�>��?Ő�D�q�Vf�7�H�)h��,21@�`{$�s�"w�i;�R��7i%K5A� mۄk���Cm��j�� �e.��ʶK�(A71o[����Dۂ�U�\^H�|��,���[Vv0�.U���*�O��N7S��Y��}j�����_G�'�@��$w2��"`h����P�a4�����4��߼(Xۺװ����l�P	4fn������'��/YȘ9{32����(��(Q���C n~r֬��$�ǹ�C���/9�ٛ�,+w�w�
��?�+J�x�v�d��怗��1��ZB��G�+�@T�f��z�����;����[��Q.n������%��p[-5z�>�����a=`A:b�ux�t�M��O�D��le�C:�z��e]���Fe�zy��Sq�1&&\�L�_=�ڪX�H~�Jנ`�b{3�K�qZ�4f_H�.1��0r�ö6�+�r�����3�Х�1�CYO>V9g�܃�����d֘���='�Q���2��S�p�h�:j��<:�Zb~UI=���b�o��-]0(ኞ&��m�c΀�O)A�uL ��l�jzYŧɹR�W��_�KB���dY�6�I�7�ו((���m�49�n��)s�XI�,j$v�@t���&�a6��O��Z[m�/\ܛ�ݵ����(����ndzD�6@3����,V�(�`�����"xL�ځ�:&�ϫ���~�A|h���t��"A��.�+u�����C��J�u�?�0/�uN=tJ	Ǆ�J���G�
���/��S�>�H
�N�+%+��ؽ��m�����<=>x��fg)��}b�����X�mN�T�ʻʯO���K���y\� ��.W�0!�\~�[���n�th�4^��[��%j�i�ĖX������ QNm�UL�5�
%��v�z#��AA�$�)%��̠,�4bH�����7������j��`¨�=0�ʖ�I�8���=���TZu�6f�Vp&��w�}X���!m��{�t떕p>����,w�y`L�3k���ޓ,21�z�m��^��'�ۍ�0k���t2P�V��(�`M�^[�6t����qu�(���k����Q*I�B��Q���/4&<�ʖ��3��bu�EØ�m�HESk��,T�)y"�F�A�d:mY�r�B\a�z��h�F��͒��q�Ň���y��$�9A���������ax��6
U*<=��M|����'Qᦣ���.�B���ͯ�_7�����H�㚹�:�xy�E,�7�֦�T����� �WA0���#��9�1$�A��n��2C��<5o	X��(Q�	vG_�\�t�5�އ#u��J�$�&T4����D���GLzRAI��6���1XASn���r}��Y��?�ڙ��@��x�/�[M{A�#ľ[�ޭ*[Nx�8G����6[�8�{�	�E��T���VXϕ��P��P,���ޕH6	f�����=\������@���I� C���VxQ���de���v^>b�mjVD�:1)m���Do�hV�{�#y��:cK�QIÕh/����z�P>⫴o�4�O�&He	]lNF/d��m��;+�恡���_sj�	�v����o��l��/�&����_w*%��:��E;��vK�{��n����.���[<U�W�߂1�:�Ff�D��Ɣ�4�?�������Yx񉋙[Y�s-Z��꼌JH�E����mt��`b��媶|��K��+9V�0J�� A0>��O��Vk�qv5bI٘�#�w���t���糮Z&��`f��#�\ج���)ӄ�i��Ƥ�zgV�5o�U��ΐS�u}N�#�� �O���nw�0}.�q�Z�8V�P�s*��̟������V��8��2(ej��������� �U���o�N�|�m.k=`(H��6�6u����#x���w��Os���H��uA�zf4�z]�E5T�
�4�H� ?:�I�)�ޔ���JEO����NV���r[</���d��)�%5��l�+�#H�srED�/���0-��+�%���.)��q�m�S��96���"�"IXZl4\���q9�l�88%��D4cV>M]zA�f(:w<ur�n����HvJ��Q�N;]�$ck��a.:ù摳5�1�&��k(�"�X�b��%����x�/a_����&4J��X�;7�xo�<��l�D�-傁Ą�G��	�z� ,��P� '�$H��"Q�,s��tJ`-������(끓��Usk����#�S˛pJl�s!Y�Q�5��d�=��h>.5�f=��x�E8��8ǈ���%o�MS�����c\��g���m{�Nq��b��J����Бl롘�n��d:���}3���G�rN�4��(.�W�Xs�O�/W���������g*��Q���@f����Q��K�,�G�VتLJ�#pv�&^>8�p�J��Vñ��x�8]�D΄�&V��2��M�=Ĥ�W��e�QAd�I)
�=�^a�Χ/��������N��R�Tˆ�2�d�y�����ŷ>1��Rb�t��f��!'�hٯB�΅pMj��_Hc�1�y���Su�㫟�! �v��뢷�r\�wZ2=s6W���U8(&�C�H�F�������I/焪�9�����j����(e2Պ�+��i%�+8��u��i�3�_�&�iE�z�3�WV	�^��xZgoT�e�R�S��� ��~�B3޺�����LM���h�Z*��@��+�Rɏ��n�����8D�0��>�.�}�)�zi�	��;t�&;����+@���Gȕ=N��(�������;�{\��x���ѼwN�-�A�?n)�C�!(o'���Nf٘�k��%Lhp��mI:Ǥ����g����ə�8g��%�iま�%4>+U�5͗=<���ާ� ?�@c�a�'���fE�襈��>���؀��ü��6]� ���[�"�<�oP�	w��á��k>�#�rZ$6W��;�Xvi�m�?�%t�px�O�ض�*2��[��S��@�}����R�9-��3	%	�=�5�T�Q�{��-Z�^�����~'�D�����Ң<�	zf�	p�U!�i�7�8r�.�i���9:��%�u�X}����ϓw���/iX����Q���=#�?"ɑ)����^e�C�x�;�j�FKʤP��Gb���T^+�y�$�wU���w8�+������� ��ᘓt�T��⺧Q|+�AV��v����S�	�F��-G��ґk>��~cց"z�%��.,�@m@?����g˪�'A(�ِ��~�x9���0	�:�GB�WC�܂bW��%2�8u������}q���r�3'���وw�����v
��:���ۅ�-���x�B����2Cmy��$~��W��\rk�	ۮt&�w�|کZ�vZ-E3��%A�HExxd�4^oh��b�k���+p��r�*�	<*�M���.�$����L��n�%�@�����t���3�� ���=�S�h+�8�s�@H��eL�'	j�=��Ə^K�>Qd3\�c�b���?�MYV�
�Nc���6�2`�{�!��`a|�ۂ9�����������o1���٘f��O�$E�OE=��fD�G/��ɪRP���U?>��g�l��|n�s���[����
��R@e^P�����!)%)��M�^��}Z�L?n�@���FQ_~�RZʎ�uT8pu�+2�R���(Dc����?Q;՘%��HU��o�z�P3����[.�ȑ�/�wl��RZ�;E�����1�n�g)�[��'jK��z�YL��D|��%�K�P��v�X̮���R�F�x�� "{.{G�Ԭ �y�qE|�>���}���c�~qzA$+�*{[n|��s�*YG;g�˄��	�2O:�0:3�o�E����};T��`J�*��m�}n���e��њF�g�#˦�Syq=�|o�H���s�����q@F.��e��S��2]C�e`�VEis/��C[�8eI�k��:veZ�Cbw	4DC���� 0i4D��2I������I}}b��d���S��Y؏"k2+ʞ5P]}z8�B�Y!�!�tK�ȥ�$�p���`��P0ʿ#���G�ߚ�l���G���{�n9��"TMF�JyS=h5�-Uo��&9�����%ڍY{�l���5Ѿߵ����=�[�>�u�K����,����e��?MN�(5:0����k�ə=�R5�ۑk�лZ�N�M� �Z�>q8��bN�S���)
�@�}��d�(�Pŧ�ʬH9d�������h���k���Z������s��Kb|E$�Aw�H�8p�Y���Ȧ���+�v;ߤ�Y�vI��1�v6���w���δ$�9����6��Ύ`_�{�/:J��J�kBG$��3z���b��M�o�� +̈́��z°sp��yL�_f�^ 9T�%Q�:�bTb�:D�J�;��DC>���y0����xg�Ǔ���gZ���`�|wC!d�Yr��3��Ŀ;�#v`��K��z0�1ۿq�(,�����ݔ���|';��Џ�9"yDr.W��Q�����w@���n�$2�#l�n�������c�"?�j'�b�ı5)~+E�4tot���/o)�-�H�9�0|��g��	^�u ���a�$����g?i8�r,i�����Q�P�6(<������I�1nӧ��(�
9����iމx�1+iV�������e�h�@4x�/uw'n�ߍ�|J�'��91��A����̃�,7p8���2�׷h��>L��J����fs��̾lݲfU��D{@��oi�~h���*��H��<�M���vH9�8���_\�ѵYF}c9���v>l�zZiP�zbm(p���΅��љ0+���D���E����0M���	}�ێ��f��q�iLD4%O�y�d�h�{��|?ON�5��g˅��,�ĒVH�"е9&�J��?�?ҖᒲT۰��E��f�R��(i=ms'Y�Ii�=Jˢ���űr�fS����?�������$n�q9o�Q��������Nq�*��gq?��#O�jzF�o�n�k�MH� ��Be���|L��g.��W����n�7@�s[F���o5����ؽ%�G��Ѹ�r"����;W��CJ�M��xL�+a���k�����'ړ��6%�L�9� ԅs�$u*)k����>{Jܺ����eg-{F�;���KYk+;E�	�f�c�iy�<%�DP$Go �˥���-Ջ{�|Y���zL�(�LR�p5�J2�1艇wC�i�^�s�C�Ӵ��Q���c}[o�;�)ت�Ye0�9�I����ǔ��Ǔ�� e���'���H'Ra��fW"@�=İ���r�ꌕ+2,�}�M�c�Ӹ8CSb��5����B���G���ǵNe8�υo,�(�q�'�����su�8MM�7$�B� ^�<:�.�j9J�A��wZHU/��G?U`��ݎ�Vl���5�%���Y4|((�z��ͭ�6����K��6bXq>!�c'��W�qn�ɡ��/�(�c�@��2ö*��V�����+�D����;��R�k�^�7�SL;]�鰈y�a� ��y�&"ضA��S8~��]�|��C+�B�a��?E22_����� ����<�D�*��V5a �G�9���[Z����}�PA+GM�����rD�\ҍz3��!��* Kt�����^����MR/����?rxJV[\��$��`ŕx%㤫�/@�K����4	�G��oqq��*Q�����l�nc�pe*aY��_H㪾F㩘_��'�O��-�y�d'�j���#Cl�Uǥ�`?{h�jpȰ`�iC�~�~�ߍ.�%s�$��	q|Q2c�'>��`��V)�������!�k�T�'e��Ak��L���'hк�}��C�r�J��`L���2�R�h�)˼&'7)a�CQ󿌃�>q��q4m�n���1*v��H/X���T�%��&�޸�f�@� 	���Q�������b�������<J�;I>�����E`���z���P�N$���`�y7�=�7y���4i�n��#u=�W�G�į؝d% �\�qi�� �I��km�� ����F��GV,4�s;�-�W`*�n����⠿�U�~�	q�}�C5W��=G�J�m��۞���@��<Κ���Qe����39U�1�:󠗽�o��qD�@���W�.�l��|�"�&�{G�估�ј�F�����a(�f�b����O��F�� �8S't,2��8�� ���O��1<a�,��QDA�Џ?+�Hӯگ�2�Mx\�,üK#��zY=���3V��y����Έ�П�#D���c-��j��(Ɨ���[��oҵ�#9g�����E����}��i;�j�[����f1�`��|�Y�h����{=���	tPROX�yK�7[�G�ٸ���;b/XYh+2��v���mϲ�:Y����3s�D@�Ng.�ұ� �����.69���rfzן��߫$;-��9������:ö��7���T$�]�Kb���Q
�\�y5c�J��/%�q&&��	S���^��ڕ�3�:| �:ר�qCG
 9�^f�CE[��r`�XT�ŐD�fB8�t�+��a���d�J-#����'��9SjQ�qP|�8�r�u�(���*�9`w
���c.��}����f�`�H+=
f)3cI�%lE���̣ii��Q،;@i6-�(�G���w}I�WT�����F!7T�H¬������� �A\(���Oe#��{���#I�*��sd}W|6ܢR�*u#���s���.z�]�"�t2A� ���%����0i܌��;�P��R�Dn���&׈|B���I.&�Hf�{0��ۆ�s,���!�w6𕭧����AC�=7�Pb_c�6�57�����x��\Ô/?��)��B],M�~�h+�F��RoQ�s�'5��	/��9D�Oe_$��u�6���ܾ,�\���,Lew>�z(�Į��X�d@���!q�M�L��x�3|�B&�����Wc�� K�����@3���a�8P��zg��I�p�Մ�OݹEPd3k�+"F�^X#���zVsҲa�Z�.fK��6ɣ��:��zw�� �n,���o5���uO@YTP�&$�L�$�@, i6���UwF�`���b�q�������/D����2�76��Ș���pV�Zh8Z�%�N�D봬�ɩI ~��"��]�5#�/N�������9�C�C�*�����oq	>�xء,p�X�c�i<5@�̆��Ż�a��X* �O��~K1+=��6�FЯe�h��`�R���Ƀڤ��	�Z��.f]m�	:R�jR;�iS|Q���D���Q(l�����5�f�����ﮩ	�d���#X��5׆5y�ͱ�=i�>���7͝]/ޞf��3�G��<�����y�*Í���ȱR�<��҉Њ p�La��.��eѿ��/�ɗ���{9��k*��⑐��ڂ)��D��c_���y�֔FKQ���"?�u���,�ńґ�e%�V�FVBAaf�W{��eRIۗ��qZ�F&*��1�@��<�܌��Tq7( ���;݅S�#V�Z��J��w"�>L�(<i~uYw�3���:��F���|�����o�h�J�'�şg��}:M!n �����'2ܖ%��-�?�W����}����%eY&�"n���w��P~��[��/�{߄�f�#�UZX�`�W�s��(z��	���̋x$����^�.�/&^,��T�[��k�Z�w���Y�M����@��p8�t�Wx��5|e��^tyxbۖ4{�H<�6��Fa�< ��S�a?x�PGY�Pvʌ!��e�o������&��\xsM�1ҳ]�j�7)���)�Z9� ��`s�o�\h�`M����/)�9b���&�.�qP�)��L��\����,��d���Э��4"ln���-��8f��gP;'y�B�ZB8"2� ����9�T�
~6�����;5�6�ėM7���W�nM5~�4�4>阽�Q��AX"�$u�	��^gHt^۷rA�u�-Z�-��OJ55�X�m���	�B�հN�`�������[�y�e�d���u �h)�C���R��8$��\�˵��>�/�"Im(�ܯ�����j��\��,铎���xi�9h�z����z}�呍���6�މIl����N��"E�XG�����O4� ����d�'$C�h����/���6j20�c��i?�2� ���.���R�J������aSE���b�R�-F)�=�~Bg��?���N�7~2B����G�O��=���D�agsc,�!ڢ�����ځk���u���p_��\�6��x�;/QI6�,�Bu�1�iz���b9?��=��%�6鉲���R7�UB3���^��ʷ�Ns2�/�A�،���W���"�y�^��@��7�
w0�&JO��'�������{���`t�@�];E�&	8x���'0�n��֧fj�O+�V����u�V�f�����.�ep|ST%�k�����]���C���-���j\w+cy��5�4	l�$�<O�������+FH�����n/��9���R��j8�j$�!08�#`}�"TI�����a��°����V���<>��~�E�f���f�36�xS	/��8g5��A��Ļ�n�����/��'�/9g��` USb�?e��3�����e�B'��"̜�����V���{�E�	�h M!�� ���~�86�X-Z>pY�-o�"H��d��PI�f��.�����\�^��VJ
$������� �N�c�r��})���z+��/{����ѧ� H���Y���2о���Y��A��C�7�/R�٘�]��+��b�B�	���u�02j^����~tv]�/�h�$��r�D:N ��[��-ȿ^�:X�bh&7��f i����R�ٱ���s29�k��ic�=~��t�H�})~r>���)Wf�&�A�^7�A
3�'��З�h�]�ZUGF؊�0�ۜ�G ~��gֿ	�NO֔��Jw���,
��e�M�r����R�)�9g.8C̀.�Օ�v	� _��-��y��� 4u�|��A��*y3������e\~��ȴ���9e�q�^y������� t7�!$%��p�Fh��4F�����LL��wY�*\JZ�S4�+��W�������B\2p&�/wkշf�ն����Fg* �˂zT~�9���Qs��t�$�Q��F�:��=&���B���ÿ�~�qT,]M�z�W�g���6�w�%��^H%��p�@����*h4Sr]��p�bd@e�T�,�	�$�z�ݶLB�J�I|�M�{&X\j�&� ��U����c���[H��{R�������#�ڸ�3������	+r=0������3��?�{r:�Ĭ�9�t6�*��+5�d�U&�l��!�-�V(�Āΐ�Ӹ�z]�?�K��H��4;�74�Nb�"k �s�7)�F&�~�?^�<e��[��{1	Ĕϛ�nf@u��#t�}Ạ�\����܃�M�A*e���8�
��
�u�}�WHz�Mﻖ,�+��� }/Tq ��]�d(,���8˪�c�PE���J/j�|J3Z�Ͼ��ôy���n���%�����(d&��;�|����z�}�J}��c��x��*��e�x��{��ܰk{��� ��K�� ��y��ѻ�u�
�^�.�t ΨL�)��p[�R�]�,�^����(���K���Ӛu��8�7��Lp�JZ1�ʥăǯw�S�v^��8�Z��4��ʡ>�s�Y����k0�	�׾���bC��A�<"qrY�Ȅs�2��]�i��S����2LG�q�����U>2�b�g��I
��u�T�LL8�A���T��J�	Swdr5����1����y��<��-o�"�nڦn�h��"$��v�;�I�lq����3�o�����"=�~�ͽ�cB�&�u0/8�[�F�D��0���3����Dͽ>S6�/g�%6��x��J^�JniΝ3۠�QR �**i��y����G\ܲ��;�FG����a����n���=�}M�U0?�w�P�H}��?���ɮ{ބKj���<�,+}/B'"D<Y|^�@" =sǬ����'&��Y�;U�ގO'd�,$F��'Z�f�X.��/ǘzR���˿;�8��E:A�G/�	��iX�)�����2�7J�O�HqM�.q ,��."vy�4j;[�ߞȪ֍�K�����UR�swZ�R�	�OT�b�"����7l�N��%����.?�� �3A�1��]3����0�����H��i�~Jg���}#_KP��]���E#��C�%����*�é���@�v��v>q+s}����9^�š5l��ߖ^�����Z���4ˏ/d ł�v��,�[d�]*��ڎTg����. ���,[+~X�ώU��Q�o�c��s?d��YA���Z&|�K>Zzr~C�ϱdo!�I�(;�J�y��RMs�9[������F!k�.�Fx��۴UB�($M'!�E8���������&Sk�=��h���G���
���ذ���J[Q1��r���h>�;���Y�q�c������8QCؿ���Ħ㜸��Y��y��)- ٠�� ��8���Ma(Q��a�\���zT��k�-\|��#f��9v�*��A(�y�H������֗�Xe����&쳶ifl����m#��?�hM�kC��P��n�,��B�(�����#	[�2�� �jw�o�f s��z�����f�pQ6.& d}5����Sp�L&�tg|�&���9�ϖ�0�{�6b�)POq[&,KQP��IG��׼�r���^$��؋��1��^������Q�+�q���D���_�m�Bv`*��p2{�cxs������i7�o�;bm%����q�����,���-�����ІsZ濏�;s�����4�1�/��;x7��c�h Sh@�R:������#a4a�|2�0����c��q�j�۴��* R�+��w]}Sw�K��c$Α��ޗ>{Ccj<M���'U��J$.�Tށ=4���Y>X��.��V��z1nE������3صY?O��l#�f�c)�KK�1n��a�Txrۺ���:�9��!�.p����}_2��'��0 j�M�k��.ڀ5t�1^���y�윔J��P���W.�JhI^j53�?��d��,�k^�Y�ݹ&Y��i�o�
�݊<����/qZ%U��'ԑ��i���CK��������N�\a=��@�,��ѳO�6���i�q�!�6Be���A�	�������/�=�}!�a-h�yO�l�%���7��&䇹A�Awud��w�rK�d�&d��#e���J�v��ӨWԲ��z�{
�ŵ+`�q�J��l��/��m!/�x�'��9(Fg W��*C����=�P���2is#�rCDC�*{Z�1FdNT8�n�6%s4�v�I,_Z�M��B[����ɛT���u;��H孬��a�1:���i�!7�"T�ؗI�.����Bv��&;y70�A.U�����ۧ`���tЅL����4�B���Da�ӝYP����n��[�Ңd&��4�_e�z��`�������Қ"��׸V.�U��I��ҫ�a��I�ĭ2­1CR<��6uBC���5}�6wC�Gۤ���/�Tc/�Y��]�#��"������'��jp�8���AǵT���[�$Z�9�қs=��$������i\}Q��2�U���z��x�f��=�',����'�&i�.�6���߀�x���C<�068�*K���C�pp���yo��ی��PTL�_�"A֚�7�HyÛ|`"TZ��?k�h������0��o��a,������#� X��\�D{8>a�K4�Rװ?&`�90����|T�kh�\�����;�v�?3����J$T��1<2!�V����{HnA�|uϞ�~�>���q�&/���������>؆�F&NT2"�����|v�J���++�����+,;�8)6><�R��Eb�1�@������B�`O�C4���ɸ��M��`Y�6��n(fL��t�^�ظD�޶��:�2�5W�c�1���EmU��Xn�2=ݪ4V#i�9OS��^y��>��KӬ:j�N�B��@H�`G�PJ9�)�6����`rp���¤�*�ú���R���9(�'jn�O�
ot��-���G�o�h��-�Z.�~
#���`#��I���z�������6��=ۗ<hFpQFR���������)�	�AXN�^b�z���âx�	4A�HIۆi����XA۫�\fJ�����놸�(�%!}�+�i�JE�3��d����t6��OgV��l �&O==�e%��Vp�j81W�FHU���^�hfFǑ��.��7@詊�{'��1]�v�@��}�����޷'�.u�[ ���wZ@�����L�!G�1D��Y��P@���`���9pZ�d��R��/�7<�(��fgX��7"Wm]!�|��$�r8��U �m�h��/����ye+e�I�!t'�s�@�3�
N�{C�#˞�va�o1�,��,��2Mٻ���K�O��&'�gm��S�,n^����T�����m`��[�y6�*�������4+�Z=O%��|����:��δ�C�r ,ۥ��"�)���#�*冐����U@_�����C����k`��������Yza�)���5-�ӫ�	��d����HL��IT�˔��q��Ϙ����m�-�h5��;L1q,�1��K41H��/��'�74ÂY������X���s��h�YZS�S�?n\�׆`<S"IH6�[Bʜ��!s�����[��^��FN����.�3���r�J{�D�|>��<qiN�>sƋ|�1N^7B���?>O'^�L+��#���V�Yad.0�1�k�z˲-�G(Y#H�:�QY�LT�m.����V��s�z��`�����O��N��Kyd2h������H~&��4?k�Hr���޵��5�=�Q�႒�W�[��&����ũ�A<Uʒ��ț�Һ{�$Tv>���c�f@s5�a���sD��R�c�^s\�����AW��(��-��+@���� ���{[������suL��P��S��7ye)�i�ٶ��
?�G��ҙ(�Mu馁��J���:Cy�rA���_⑎i��K�����n5�Ou���;P~s�ČKS�gy��fu�H��/���xL�y1l)^�O�{X�/!�'�z��僃C���|�&|%�1��m%@1�e�Y�[�6�� F����x@K�
aIF`�`HI��g�b�5��x��/���щ�K{�_��)$ރo�D�)u��,��ķ;v]��
��L���} M:/���xP�q�i6B��n�upPC>"ʮ�
�sg�d~�XK%�Vjn4� �,�,٠��i	"��gZ%Ь]��i	��4S�b������-YS�e�yɚ��i���M_��GZ�ɸ������)T��-�l�tVM�Ŧ���X�X`o����?X��!���m&:u�"���K�j������=x���=IM�>r��4>(<�>��w�´��p��$Jr���p;�������0St�]��*��Y�g�c�Sa�i����d�C@GV�$�`	�WΈP�K_4��!:���h�_.�d�2Zd��^����Y�\�G��.k�B�>�d�z�l����:�Hg�o����_K-~�$��1��M�^��(�ZNj��:����V��*Lǵې�V������Bn���{�k.����]osҿ�pk�c?r��=.p���sUq:�v��0N�ʔ�"s	��p��3B@���b���MS/h0�H��s���s�e<_�<}n��NG�*�E���!Mm�b���Z�X|�<g�'s#�-3x5��2�g[΂bI׹K$����|C�aa��\Pm\�1��]jR��#�E펤}�������x��]����/`uvW�w�L�)CvwT�,�tS2���#����E�@=6e:1Y�Q	�?��i�sC��(��5�rD*o���Q#�iynkJ��;^�	+�%FL�B���4�Pmi�� &�²�>�a�u����7�a\����+"�l�!���XgYzE:"�X(vS��0�WXdȶN�D�	R.3Aw�i�B�b{ϳ��Wyj��r�u�t�G�v9�Qx2�^Xy4]�\]T�ɡ@
\;��.��s���ǅ�b�Q[�|��U��v��zn�zNG�`������Igk����0�e�r��3Tx�",��
.�u9;Z`�yc����h����c
jػL�Fb/�Y

�.z��,�Q���L	�*Hd�U���uOq����me߯Ι��rѶ��"�Q�y�W�%tϙ�BPVR��/.Pe�!����,�����d�J�Q���]���ߕ��<�	K/*���pS�-8vm�1}����jZ(U+j	��F�xZe�n���)�E� ]^~D����+��������+93�t{�T,ݢ<|h\�}����L��Z-5�;��[�e�p�'!UC�c���f�ea�~�L&g��1lO��".}�S�=�>�}/��Н@x�&���!�)Yq���"�c�;T�I����X�d�O�Z�K�R�Kqҹ/f�US��<C�����I�L����j�e�H6���/mYd=��֦�tnd�`1 ��i٧z����ֽK�����Ë�/}8���U����G�Q���%�6̝�5����٘�΀D��k�A�e~م�.�䳝�#>��L6f�k$�G�>ט�D����wo���_{�ɡ����^����iNq�����(�@��З����7�kY��J �g�	lӈ���,����?�G�K*7N� tR��x%��x�5��nSW��0�;��h��-�D�dϷl��X��}pU(�ܭ6B�"o��/��.��%�K*-������)E��D�-�{7��RqϽ��RΜ�϶��rOF�Z+���FLn��v_u-^c"�nk���8Auc���O4��f�;G���K�dv��Y��L
6��1�*�aVy7��}!M�N�,0A�s�0r�����I�/�W�%��c��#I�p�i�(�c�Xt	|�a1����/��\�(:����]�@⺌�$%i���b���R�f���~�!%Y����~��7�6N��r�לu3��϶]Yx���ֳ��}�>oW^lw�LL)i�c�7D,�s譌��]�E����D���z>qn�ɉì��/9dC(7Wk��ZٻCR ?�ҵP{)�����C
wp{a2� D\!�t#
����b�3�����po��t��>L�ȃ�����\L�~�e�):n��:&s���o�����~�H���g����rdQ;�`phf �����c�0�� ��!֤M�Aha<�� +n��u�	V��')����,2W23�\:�l�0`�P��"�����}��#5���Q�8JLg��g�W^�q���y� y�X;���y���3*��% 2�}���RP���u��w����>ZmRq�'���#Z�cJ
�Y|��������bư����#{�%���A��".�o�3�v�-=���g$b������<="�h���9Cė#����]�:JPRu�/̍s��Q�2����+ɦ}�ħ�J�o�͐?��I��#16.�a�Cf�ܩS _��oO��V$���>�dƺ�[*{KG�+����ɲ���J�15N�)S2 ��{�� ���C�7��ۖ��>PL}��=��Dӭ� o���6�s�j:�/<l����a�!�}�Y��L�L��J��3T�� �|䉉q�-��H���v3x?Bk�K�#�SP�������r���J�H!����zKW�h�؇a����U�6�r��	�@9�����b�&#�5�@��n�^+�7��5���Zя�Q,5�<�ft��{F����-�����a���46!+�e�Aވ'�d���%������^e�D���&C��F�U.���CY�P�c�{�fƸ��W���s�=iat}��:� &-��rYa�C��[�1/��%V6�3_�
H�M��j`�	�~R�\���7�)�bzI�JnƯ7�\rч9h0��;�z��%-W�Z5�.�V�$���.{��G�K&����8M�.�N���x�S��M��a��_�8oTd�:�)9V�ot�M\�ߍx��=1P?E,2M�c�*]a�$ѡP\aS���_|�)���@�Z��x?X�����4e6��6|˾���\q�������!Jn:^��i�9g)"ww�����p���y�o�1�	�����2H�,{�L�wq�TMXbJ��iQ�iͲi_���=u!Ew�G4�X�n
pӳ�k����d��)3��]�H_��lM墚7�w~i�qVR��o�:٢��1��P�7H�}�FIb���V[ ���x��Z�G�m��O_zp��r�W�NY���zt8�s�0:/u�\�+��1H���
��,�c"�՘�o3����N!l�,.��xȒ1W����/Lg�{���8kr��Oͪ��ۅ�)�*���f)�*��B�`���eK�p	�������!y���I�5�Y�����l.��m�I��|x�DF�:�\R�7Ve �r5�L�6����K�$�A��Y�h�E��XOw��� 
�C�卷�^��Ë❝��o{a�n�\����gU��Dn�pЧB��z��JF��Q��A��hu�2��:���1��J��V����x�%� �\F!��xO�:��=g�Խ*�,u�K�3���亜�S�X?���0�� 
Uv>�א��),b>��@$��m���V:�� T���0r���2Eў��*a�dJЪL� lU��1�S�9�����0��1ܒ�NK�i}����:-����Yg,����4�_�~L1�+���3!A��T�\�O�\&�gx��N�)�Mq�0�6/�m$6�(��~d�9g	_/��'���TV��Z�<�}�И�uV	Nݮ��$��,_��"K*�>�+����B�z��T���Uto��q��n�=�=>�x�BQ'?J$�:�He��.����*���V�}Q{�	�Ȝ��Y��٨CP��Rn���g���T�D4ﶈ���Cg*���v�;�p$��5�cڠG�j��J��B�kjYa�%s�2šs��le!��bgn����~�ť��@��]9Z.�p�l]��a�0y��]���'"~�a��Jv�� �J;itBv�_ں���=1
�V!����A �_V�׳h]s�O�QT0��sX�_M�e�]����+�#/�~�tWO������x(;ۍ���g4E�đ��̻M*SE\+�Q��&{���*6�<�#l��Yj���QHT(�Jg�m��ޔ�=�V��Z@l�{��-]������k	>��z��3���.�q���H��D0;H�H�
�A�D�y��?��P����=�����;'.t(��`�N�l!��?�oWz��E��I��H���n>��$�� kbs}�b�iJ�R���;C��0�4���� ��k�
��_���D�� >d;-�?���RhZ�$P���W�Xgl���ǔL����Pp��s�yd�IR��h����-�7WZcF��1���:8�Z���!qV�M���������oum�%�*f`�.5I�@Kp��)D������U+-߸ 83"8�F�߹]&%
Ρ �Ʉ������ k M膆���O��
/�h��!�V��K�n=����Vڊ���2�B��Q�?;z��@����un�_�8]�)���k�uI0�Z�=�{��� �Z�y�V��!���h���?/Eߝ�]�N���PP��â�er� �x����Qsy}���{$g�'j�>�+߅l`���D�#�snrOG+F�<��L�b�J�r������g�Sڳ�-4j&P�L���$��8I\�s5�w�<�����ƭ��L\��|=�!\��%��^�k�d��P�!#~k���3�M��]�g�%;�=�`S�c� 2��z~k:���s)+=6ʒd�����W�'�m��,L��ɪnL6�A�3��N�z0����\�"9���o�j��S�$�q��s�'(�Ʀ�RFS\q����	� �C�6�m���F�
��mӵ��ɸW2��� e591iO�0���A�g�`Q�K*�P���:#���7��U]��u����ը�����E$aל�?8(R��a��'���z���3�}����n! S���[б<��]i���~]1x��f// ������	�M��3���Ě��]g�ă�h����`�k]ɫd�V��Yo�%�������ϓTe����^����F�Ki��xP�����R�V�NڰOtt�A�EbѲ��|�17�����j��8�k��m�F�r*�̮��tJ�Q�K
����LVUԼy!����q�����u	HV�����U�sSp!v�e*�4�\S��Q���b�4�����m��\�&@^�М���y��r'�lb#����@v/U�Ȝ�U~.��<N_/�7��꣢�H�h\8��u��z��]_�a�����<�����P���s8k���	�D��n �2�/��$�r!\�ۯ?�j+�(�C�g9]i;�iM'��c��M��|����D�2Uʃ*���CWD -�D^ ��Ƭ�Z!�~����Tf� ���{.��UO����Hy=#�/�&�Q�r�?�k����~��g/��8w\��;�.���W^v�s���H7�b���5AA5�-HSĦ�(7�{���ȼ#�V|�
���2���e��iD�I�iSB�_����#�
�����N?́k��^��-b���\m�b�<�c?L��_B̹�q�N�g��۟���M,Ig��mv�� !@��-��ܣH�]Ƕ-�0,�� ��|D8FL�?S5��hlHI�".�eN�ៈ��@���0���El	j��/�̹�UuؾgⓅZ7����;M�@Gjey �_�XnP ��Dm��j�;�&�dH�Z����9á�%�,�n�.���=�1��Z�� �
�d�9��?�j�+a#�G""f9�4��>-�M�0r8_�!f��O,J�D��'�� ��{�@�&q�(������,��,�81�A �i�?�U��,P�� 'R�_�����p��]y����L���8/�+%��Me�
�;h�
L'����M�)`�#p�×��Fs��nٝ偩K���ݾk�%KB��Gu�I�ъz�#KqR0 >ay��n�c5χUR�q����X5C�d�a(wz�5�y��j�xs��֯p<���U^3+|q�P�e(���&�	d��a`�G^�"�4Ƶ=џ�s��_����O��l����t���0�q*W��r�f�*�o�PFc�X�c {
�B�O|�}_,����5Xb�6�4�/�W�RkÑ_�52�ah�l����N~�5�����������-�����5K���u�W���ڮz���_{R����_�Y2�b�N����'79Tb(TO?p[Ja������R����5R��+�:��Ί����"/�x2�.�S�����׮�4P��a$��$���7���D�~���4?|��f�e�u�Ѱo��V<�>�Am��к���RT���z���7(�=�:�-i�V��;І�P�M���G�y\x� @�-Z�Ά��|���Ǉ��Uy��,e&Ⱦ��.����"Ytv[�+@IZ�_Ib̔���]���w#R�6c��<��&�	���)@Hd3i�y7a.P1���l#���Nq�s�C�g#�}�%p�<��67�Dʹ��)�k��(�E�9�4�;�R����|�@d���sR>���x���*�ؤe�p�~(�g ySF�������)'�݄C�E~��Zz&�q��`�����5	�}�Z\]c��+[�6n�`1�k;zEb��V7�m�J0��~zy����Y�J㫢�e��1K�.\����I�h]گ�U_�*�Cp���:jr:R�8�s�}��J��v{�ͱ�8Z�C���c=����8����d?q�����R4��`�+'ʇS@�����Ӫ�����z	Ʊh�����I��g�5A Y��yu�_5�͐�a�5�rv3�K	�<L�"q�|����+>)��a�7j����h�AHOUS!��)�EN̎������T�}w�g���b+��� N�E�L65�0U�:T5{��tl��)�;�J�)�d���-^��kne]^��T���	�����fg��kϣ^�ɞPp�g&X���E�E��E�5
��VJx�EpF1�t��W����C�[����0�:&����i#%�9*���b���瘧�/�o��
��s���ޥ��L�
^�j[��v�
7X����($'�"��s�Ӿ�7�P�&,]���T �7�Ӆ�ȳ���$Z H,�e@�h����v�]���K�Ʀ#,��ޑ3�����a" 2/��w�.���]�^)1�I����A;`k�[��W�32���u�8����:�=��ق9��V���Wj���`� D9h�N���Whd�m�t�ƞ]�	ws�|������g�^�~��@�^��(���4�u$��n��W�r����X���/�Vo�o.�0!�1$�vn��)�t�V��~��h+a3z��ޚ�/�`6�6	&bA�Ϻk��6�m�q]�5R[U�����z�.�H�3LT�+��3��,��Jv6����ڪ�Qb#�JK,�K7��l��1���'���0�o�n������*a}�����u��6�|��H�����Jc�ö����=���ݗ�&���l���s�B�����JW���й��w�tE%tv^�n�!��jGK)�ovZ߮)O�O��f��/x-~��v���ڴ8����В3��.d�J'r�Di��G��������S#��d �>�{ю?���B%��I0BѸ<��
��} �.��m�~,�y*����G����3%��zyk�� �n��Z�ZꉬV�?q�`��e|��X%�a?^YM�=�)a��T�ʅ�ܿj
(u�F������y��.���'
�`��5��f�vZ%��̖͵����$�ur����3>�&p�f��n�@N�dE�CE]a<����[��7���l�K��\~6nP�������q��i����s��]%X�ąy�`L�nJF�)��d0R�7�y�ϵ>w��K��iJQxVm����:[��Np�M�=m�'#�g���Ll����f�P�z�6u��H�ne��?D�+d$m�=��[��@���>�_����%�p��AEoV��k�X��|8ݣ�"G��Y��</��n��i���U�=���7S��r&tT��|mM���ɽ��4�A���v���T���U� gr	E����z6Q�V��#�h���A���q�� ��q)MJ��~NCXF��w�9@Ar�!�S
�|�M1�n8��2����p�lh_4��Q�=�c�R�*c/�r�MҤ�B��v�V�-W�&�G[a��d�(�RV��#�d��
������JȟQK�ь%#�O}�w��^��<	%��Qi���e�0��owsp���8��Cr!y�eb3h�I��>�����zJ|�]��v�S���
2Y)���bt�rd�ZQ4�XB-ׇ��!,��-[~��Sz�,��0fE�M�d�"�i����~���B�"|̐�n�Z?�%�}.3�|��OE봃�H+���鞓X79�<�o&�78x�|P�%�D0
bh��� ��P�}�s�D�n����r�+�[�)��%+P�~II�Y�!��a�d�̢�GQ��M�1��Љ2���a��l�;�I:��(�S��i������=B-H�Z�
����>*ҎQ�85�1s^p���d�nkU+�yF���W�U����Q��~(�蹖��w��N����)|�Ǐ̟$����$��PN����M ���l(���Z��&��?��^�feMaMZV���T�����YIW��Z�ťf�vh&���]� §���=����md���I �B*��
K����$���"c�ɠ�l���p����u����q�	[Q��/�����k�^\ ;f�:,��r��3�Q�zda�H�A'�&����=��a���1	6��=�@� ,�[(�Qn�=�Q��p
[�롯�<���7�	�M����Q�u����n�y���
����5��F���$�v�4Q��Iڿik+�0���(v��L�ƴ0|�:��(�Y𺭾���i6�����	%��RX���HH�Em�Le���N�O����r�rEP�����M��D����:�㊎O|�k$lS���~)�f�����C�#*Q�z�n�t�yu-����2��������UV�+SC�ꚑ|�-۽��ف�=Ah�(�y7.Q ��'�{F_�����a�v �Wu�Uc�0���|�>*�N���5
��ڐ�V�s���a��V����Ex�A�u_ؑ��Tj�v@�k�]����%`t�"+�E�1��x��::[�{&&9]��C��Η�����sz�Wq��A���?6jI�Wx�JjM^���n#E�|G][��A+Σ:�ϵ��
�m��_x<�k\�Y���{ ;b~��Qy�c̷h��Soƒ��9h}=����ԍS��­�&��$� ���{
%l��fO\(6܀�s�/�qc�g-ke��{][$�t�*���i���:���j4�W����~�G�Z۷A��SU�(6\���a�.�PKjO۫�q��Nfh��m�)��5�vZ�@���%N�X��c���GV͋ϖ���\���]�w�I��F���j�:�c����hPN���7���F��ϯ${���ď�6!L�_vX&�MU�č[c^����x5u$:��/Tj�xp��$u����rOd��Ce5N�P��͹�D�λ3�p�`VȂ6i��������u�
�DH�8+3������ Ki���s�7��[>-���b�����U�*世ȡ���>]%��Ή�{�8Dnz?��I)y��`Rߴ��Ĳ�>�	@���Ts���¿��8"��q14��/l�,���*��<�X�fp(%GA�j�����3���,N��K�	�Q�X��CA�N�����0]�g�VY�7�c�>|��b���/��J������̊��^�S��'����2$�Ӥ���$��0�!%c�Z�rΖ��ѭ�ځ�o��:x��g�ܷ���aY.fZ�S��	*�&�kܘ{#!��8�ms��I��LHHe�y���N��co��C(;�_� �#	��*0[{U��{��ǧ���i�vdΕ�*qJt��Oe�#����ttI�·�O80��Ώ�EJ�e�T�$��s�B{�HS�?�U?���$�r��=����d=�QF�p�#��$sBh��d���B!c����k��ni
T�Y���~)� �V	��|�)�i�s��t'����K)+@��� ���΀/�(ڨ����Y��C�C�S#M�u���������"���C��k����Ha�J�