-- nios_tb.vhd

-- Generated using ACDS version 13.1 162 at 2022.11.16.15:37:35

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity nios_tb is
end entity nios_tb;

architecture rtl of nios_tb is
	component nios is
		port (
			clk_clk                          : in  std_logic                    := 'X';             -- clk
			pio_0_external_connection_export : in  std_logic                    := 'X';             -- export
			pio_1_external_connection_export : in  std_logic                    := 'X';             -- export
			pio_2_external_connection_export : in  std_logic                    := 'X';             -- export
			pio_4_external_connection_export : out std_logic_vector(7 downto 0);                    -- export
			pio_5_external_connection_export : out std_logic;                                       -- export
			pio_6_external_connection_export : out std_logic;                                       -- export
			uart_0_external_connection_rxd   : in  std_logic                    := 'X';             -- rxd
			uart_0_external_connection_txd   : out std_logic;                                       -- txd
			pio_7_external_connection_export : in  std_logic_vector(7 downto 0) := (others => 'X'); -- export
			pio_8_external_connection_export : out std_logic_vector(7 downto 0);                    -- export
			pio_3_external_connection_export : in  std_logic                    := 'X'              -- export
		);
	end component nios;

	component altera_avalon_clock_source is
		generic (
			CLOCK_RATE : positive := 10;
			CLOCK_UNIT : positive := 1000000
		);
		port (
			clk : out std_logic   -- clk
		);
	end component altera_avalon_clock_source;

	component altera_conduit_bfm is
		port (
			sig_export : out std_logic_vector(0 downto 0)   -- export
		);
	end component altera_conduit_bfm;

	component altera_conduit_bfm_0002 is
		port (
			sig_export : in std_logic_vector(7 downto 0) := (others => 'X')  -- export
		);
	end component altera_conduit_bfm_0002;

	component altera_conduit_bfm_0003 is
		port (
			sig_export : in std_logic_vector(0 downto 0) := (others => 'X')  -- export
		);
	end component altera_conduit_bfm_0003;

	component altera_conduit_bfm_0004 is
		port (
			sig_rxd : out std_logic_vector(0 downto 0);                    -- rxd
			sig_txd : in  std_logic_vector(0 downto 0) := (others => 'X')  -- txd
		);
	end component altera_conduit_bfm_0004;

	component altera_conduit_bfm_0005 is
		port (
			sig_export : out std_logic_vector(7 downto 0)   -- export
		);
	end component altera_conduit_bfm_0005;

	signal nios_inst_clk_bfm_clk_clk                              : std_logic;                    -- nios_inst_clk_bfm:clk -> nios_inst:clk_clk
	signal nios_inst_pio_0_external_connection_bfm_conduit_export : std_logic_vector(0 downto 0); -- nios_inst_pio_0_external_connection_bfm:sig_export -> nios_inst:pio_0_external_connection_export
	signal nios_inst_pio_1_external_connection_bfm_conduit_export : std_logic_vector(0 downto 0); -- nios_inst_pio_1_external_connection_bfm:sig_export -> nios_inst:pio_1_external_connection_export
	signal nios_inst_pio_2_external_connection_bfm_conduit_export : std_logic_vector(0 downto 0); -- nios_inst_pio_2_external_connection_bfm:sig_export -> nios_inst:pio_2_external_connection_export
	signal nios_inst_pio_4_external_connection_export             : std_logic_vector(7 downto 0); -- nios_inst:pio_4_external_connection_export -> nios_inst_pio_4_external_connection_bfm:sig_export
	signal nios_inst_pio_5_external_connection_export             : std_logic;                    -- nios_inst:pio_5_external_connection_export -> nios_inst_pio_5_external_connection_bfm:sig_export
	signal nios_inst_pio_6_external_connection_export             : std_logic;                    -- nios_inst:pio_6_external_connection_export -> nios_inst_pio_6_external_connection_bfm:sig_export
	signal nios_inst_uart_0_external_connection_bfm_conduit_rxd   : std_logic_vector(0 downto 0); -- nios_inst_uart_0_external_connection_bfm:sig_rxd -> nios_inst:uart_0_external_connection_rxd
	signal nios_inst_uart_0_external_connection_txd               : std_logic;                    -- nios_inst:uart_0_external_connection_txd -> nios_inst_uart_0_external_connection_bfm:sig_txd
	signal nios_inst_pio_7_external_connection_bfm_conduit_export : std_logic_vector(7 downto 0); -- nios_inst_pio_7_external_connection_bfm:sig_export -> nios_inst:pio_7_external_connection_export
	signal nios_inst_pio_8_external_connection_export             : std_logic_vector(7 downto 0); -- nios_inst:pio_8_external_connection_export -> nios_inst_pio_8_external_connection_bfm:sig_export
	signal nios_inst_pio_3_external_connection_bfm_conduit_export : std_logic_vector(0 downto 0); -- nios_inst_pio_3_external_connection_bfm:sig_export -> nios_inst:pio_3_external_connection_export

begin

	nios_inst : component nios
		port map (
			clk_clk                          => nios_inst_clk_bfm_clk_clk,                                 --                        clk.clk
			pio_0_external_connection_export => nios_inst_pio_0_external_connection_bfm_conduit_export(0), --  pio_0_external_connection.export
			pio_1_external_connection_export => nios_inst_pio_1_external_connection_bfm_conduit_export(0), --  pio_1_external_connection.export
			pio_2_external_connection_export => nios_inst_pio_2_external_connection_bfm_conduit_export(0), --  pio_2_external_connection.export
			pio_4_external_connection_export => nios_inst_pio_4_external_connection_export,                --  pio_4_external_connection.export
			pio_5_external_connection_export => nios_inst_pio_5_external_connection_export,                --  pio_5_external_connection.export
			pio_6_external_connection_export => nios_inst_pio_6_external_connection_export,                --  pio_6_external_connection.export
			uart_0_external_connection_rxd   => nios_inst_uart_0_external_connection_bfm_conduit_rxd(0),   -- uart_0_external_connection.rxd
			uart_0_external_connection_txd   => nios_inst_uart_0_external_connection_txd,                  --                           .txd
			pio_7_external_connection_export => nios_inst_pio_7_external_connection_bfm_conduit_export,    --  pio_7_external_connection.export
			pio_8_external_connection_export => nios_inst_pio_8_external_connection_export,                --  pio_8_external_connection.export
			pio_3_external_connection_export => nios_inst_pio_3_external_connection_bfm_conduit_export(0)  --  pio_3_external_connection.export
		);

	nios_inst_clk_bfm : component altera_avalon_clock_source
		generic map (
			CLOCK_RATE => 50000000,
			CLOCK_UNIT => 1
		)
		port map (
			clk => nios_inst_clk_bfm_clk_clk  -- clk.clk
		);

	nios_inst_pio_0_external_connection_bfm : component altera_conduit_bfm
		port map (
			sig_export => nios_inst_pio_0_external_connection_bfm_conduit_export  -- conduit.export
		);

	nios_inst_pio_1_external_connection_bfm : component altera_conduit_bfm
		port map (
			sig_export => nios_inst_pio_1_external_connection_bfm_conduit_export  -- conduit.export
		);

	nios_inst_pio_2_external_connection_bfm : component altera_conduit_bfm
		port map (
			sig_export => nios_inst_pio_2_external_connection_bfm_conduit_export  -- conduit.export
		);

	nios_inst_pio_4_external_connection_bfm : component altera_conduit_bfm_0002
		port map (
			sig_export => nios_inst_pio_4_external_connection_export  -- conduit.export
		);

	nios_inst_pio_5_external_connection_bfm : component altera_conduit_bfm_0003
		port map (
			sig_export(0) => nios_inst_pio_5_external_connection_export  -- conduit.export
		);

	nios_inst_pio_6_external_connection_bfm : component altera_conduit_bfm_0003
		port map (
			sig_export(0) => nios_inst_pio_6_external_connection_export  -- conduit.export
		);

	nios_inst_uart_0_external_connection_bfm : component altera_conduit_bfm_0004
		port map (
			sig_rxd    => nios_inst_uart_0_external_connection_bfm_conduit_rxd, -- conduit.rxd
			sig_txd(0) => nios_inst_uart_0_external_connection_txd              --        .txd
		);

	nios_inst_pio_7_external_connection_bfm : component altera_conduit_bfm_0005
		port map (
			sig_export => nios_inst_pio_7_external_connection_bfm_conduit_export  -- conduit.export
		);

	nios_inst_pio_8_external_connection_bfm : component altera_conduit_bfm_0002
		port map (
			sig_export => nios_inst_pio_8_external_connection_export  -- conduit.export
		);

	nios_inst_pio_3_external_connection_bfm : component altera_conduit_bfm
		port map (
			sig_export => nios_inst_pio_3_external_connection_bfm_conduit_export  -- conduit.export
		);

end architecture rtl; -- of nios_tb
